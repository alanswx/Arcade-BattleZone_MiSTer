wave_lengths[0] = 16927;
wave_lengths[1] = 16942;
wave_lengths[2] = 16958;
wave_lengths[3] = 16974;
wave_lengths[4] = 16990;
wave_lengths[5] = 17006;
wave_lengths[6] = 17022;
wave_lengths[7] = 17037;
wave_lengths[8] = 17053;
wave_lengths[9] = 17069;
wave_lengths[10] = 17085;
wave_lengths[11] = 17101;
wave_lengths[12] = 17117;
wave_lengths[13] = 17133;
wave_lengths[14] = 17150;
wave_lengths[15] = 17166;
wave_lengths[16] = 17182;
wave_lengths[17] = 17198;
wave_lengths[18] = 17214;
wave_lengths[19] = 17231;
wave_lengths[20] = 17247;
wave_lengths[21] = 17263;
wave_lengths[22] = 17279;
wave_lengths[23] = 17296;
wave_lengths[24] = 17312;
wave_lengths[25] = 17329;
wave_lengths[26] = 17345;
wave_lengths[27] = 17362;
wave_lengths[28] = 17378;
wave_lengths[29] = 17395;
wave_lengths[30] = 17411;
wave_lengths[31] = 17428;
wave_lengths[32] = 17445;
wave_lengths[33] = 17461;
wave_lengths[34] = 17478;
wave_lengths[35] = 17495;
wave_lengths[36] = 17511;
wave_lengths[37] = 17528;
wave_lengths[38] = 17545;
wave_lengths[39] = 17562;
wave_lengths[40] = 17579;
wave_lengths[41] = 17596;
wave_lengths[42] = 17613;
wave_lengths[43] = 17630;
wave_lengths[44] = 17647;
wave_lengths[45] = 17664;
wave_lengths[46] = 17681;
wave_lengths[47] = 17698;
wave_lengths[48] = 17715;
wave_lengths[49] = 17732;
wave_lengths[50] = 17750;
wave_lengths[51] = 17767;
wave_lengths[52] = 17784;
wave_lengths[53] = 17802;
wave_lengths[54] = 17819;
wave_lengths[55] = 17836;
wave_lengths[56] = 17854;
wave_lengths[57] = 17871;
wave_lengths[58] = 17889;
wave_lengths[59] = 17906;
wave_lengths[60] = 17924;
wave_lengths[61] = 17941;
wave_lengths[62] = 17959;
wave_lengths[63] = 17977;
wave_lengths[64] = 17994;
wave_lengths[65] = 18012;
wave_lengths[66] = 18030;
wave_lengths[67] = 18048;
wave_lengths[68] = 18065;
wave_lengths[69] = 18083;
wave_lengths[70] = 18101;
wave_lengths[71] = 18119;
wave_lengths[72] = 18137;
wave_lengths[73] = 18155;
wave_lengths[74] = 18173;
wave_lengths[75] = 18191;
wave_lengths[76] = 18209;
wave_lengths[77] = 18228;
wave_lengths[78] = 18246;
wave_lengths[79] = 18264;
wave_lengths[80] = 18282;
wave_lengths[81] = 18301;
wave_lengths[82] = 18319;
wave_lengths[83] = 18337;
wave_lengths[84] = 18356;
wave_lengths[85] = 18374;
wave_lengths[86] = 18393;
wave_lengths[87] = 18411;
wave_lengths[88] = 18430;
wave_lengths[89] = 18448;
wave_lengths[90] = 18467;
wave_lengths[91] = 18486;
wave_lengths[92] = 18504;
wave_lengths[93] = 18523;
wave_lengths[94] = 18542;
wave_lengths[95] = 18561;
wave_lengths[96] = 18580;
wave_lengths[97] = 18599;
wave_lengths[98] = 18617;
wave_lengths[99] = 18636;
wave_lengths[100] = 18655;
wave_lengths[101] = 18675;
wave_lengths[102] = 18694;
wave_lengths[103] = 18713;
wave_lengths[104] = 18732;
wave_lengths[105] = 18751;
wave_lengths[106] = 18770;
wave_lengths[107] = 18790;
wave_lengths[108] = 18809;
wave_lengths[109] = 18828;
wave_lengths[110] = 18848;
wave_lengths[111] = 18867;
wave_lengths[112] = 18887;
wave_lengths[113] = 18906;
wave_lengths[114] = 18926;
wave_lengths[115] = 18945;
wave_lengths[116] = 18965;
wave_lengths[117] = 18985;
wave_lengths[118] = 19005;
wave_lengths[119] = 19024;
wave_lengths[120] = 19044;
wave_lengths[121] = 19064;
wave_lengths[122] = 19084;
wave_lengths[123] = 19104;
wave_lengths[124] = 19124;
wave_lengths[125] = 19144;
wave_lengths[126] = 19164;
wave_lengths[127] = 19184;
wave_lengths[128] = 19204;
wave_lengths[129] = 19225;
wave_lengths[130] = 19245;
wave_lengths[131] = 19265;
wave_lengths[132] = 19285;
wave_lengths[133] = 19306;
wave_lengths[134] = 19326;
wave_lengths[135] = 19347;
wave_lengths[136] = 19367;
wave_lengths[137] = 19388;
wave_lengths[138] = 19408;
wave_lengths[139] = 19429;
wave_lengths[140] = 19450;
wave_lengths[141] = 19470;
wave_lengths[142] = 19491;
wave_lengths[143] = 19512;
wave_lengths[144] = 19533;
wave_lengths[145] = 19554;
wave_lengths[146] = 19575;
wave_lengths[147] = 19596;
wave_lengths[148] = 19617;
wave_lengths[149] = 19638;
wave_lengths[150] = 19659;
wave_lengths[151] = 19680;
wave_lengths[152] = 19702;
wave_lengths[153] = 19723;
wave_lengths[154] = 19744;
wave_lengths[155] = 19766;
wave_lengths[156] = 19787;
wave_lengths[157] = 19809;
wave_lengths[158] = 19830;
wave_lengths[159] = 19852;
wave_lengths[160] = 19873;
wave_lengths[161] = 19895;
wave_lengths[162] = 19917;
wave_lengths[163] = 19939;
wave_lengths[164] = 19960;
wave_lengths[165] = 19982;
wave_lengths[166] = 20004;
wave_lengths[167] = 20026;
wave_lengths[168] = 20048;
wave_lengths[169] = 20070;
wave_lengths[170] = 20092;
wave_lengths[171] = 20115;
wave_lengths[172] = 20137;
wave_lengths[173] = 20159;
wave_lengths[174] = 20181;
wave_lengths[175] = 20204;
wave_lengths[176] = 20226;
wave_lengths[177] = 20249;
wave_lengths[178] = 20271;
wave_lengths[179] = 20294;
wave_lengths[180] = 20316;
wave_lengths[181] = 20339;
wave_lengths[182] = 20362;
wave_lengths[183] = 20385;
wave_lengths[184] = 20407;
wave_lengths[185] = 20430;
wave_lengths[186] = 20453;
wave_lengths[187] = 20476;
wave_lengths[188] = 20499;
wave_lengths[189] = 20523;
wave_lengths[190] = 20546;
wave_lengths[191] = 20569;
wave_lengths[192] = 20592;
wave_lengths[193] = 20616;
wave_lengths[194] = 20639;
wave_lengths[195] = 20662;
wave_lengths[196] = 20686;
wave_lengths[197] = 20709;
wave_lengths[198] = 20733;
wave_lengths[199] = 20757;
wave_lengths[200] = 20780;
wave_lengths[201] = 20804;
wave_lengths[202] = 20828;
wave_lengths[203] = 20852;
wave_lengths[204] = 20876;
wave_lengths[205] = 20900;
wave_lengths[206] = 20924;
wave_lengths[207] = 20948;
wave_lengths[208] = 20972;
wave_lengths[209] = 20997;
wave_lengths[210] = 21021;
wave_lengths[211] = 21045;
wave_lengths[212] = 21070;
wave_lengths[213] = 21094;
wave_lengths[214] = 21119;
wave_lengths[215] = 21143;
wave_lengths[216] = 21168;
wave_lengths[217] = 21193;
wave_lengths[218] = 21218;
wave_lengths[219] = 21243;
wave_lengths[220] = 21267;
wave_lengths[221] = 21292;
wave_lengths[222] = 21317;
wave_lengths[223] = 21343;
wave_lengths[224] = 21368;
wave_lengths[225] = 21393;
wave_lengths[226] = 21418;
wave_lengths[227] = 21444;
wave_lengths[228] = 21469;
wave_lengths[229] = 21495;
wave_lengths[230] = 21520;
wave_lengths[231] = 21546;
wave_lengths[232] = 21571;
wave_lengths[233] = 21597;
wave_lengths[234] = 21623;
wave_lengths[235] = 21649;
wave_lengths[236] = 21675;
wave_lengths[237] = 21701;
wave_lengths[238] = 21727;
wave_lengths[239] = 21753;
wave_lengths[240] = 21779;
wave_lengths[241] = 21805;
wave_lengths[242] = 21832;
wave_lengths[243] = 21858;
wave_lengths[244] = 21885;
wave_lengths[245] = 21911;
wave_lengths[246] = 21938;
wave_lengths[247] = 21965;
wave_lengths[248] = 21991;
wave_lengths[249] = 22018;
wave_lengths[250] = 22045;
wave_lengths[251] = 22072;
wave_lengths[252] = 22099;
wave_lengths[253] = 22126;
wave_lengths[254] = 22153;
wave_lengths[255] = 22181;
