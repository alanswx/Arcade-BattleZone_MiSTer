jegor@Jegor-Laptop.390397:1613475082