squeal_samples[0]=28998;
squeal_samples[1]=31377;
squeal_samples[2]=33654;
squeal_samples[3]=35834;
squeal_samples[4]=37910;
squeal_samples[5]=39903;
squeal_samples[6]=41799;
squeal_samples[7]=43615;
squeal_samples[8]=45354;
squeal_samples[9]=46905;
squeal_samples[10]=48403;
squeal_samples[11]=49919;
squeal_samples[12]=50103;
squeal_samples[13]=45584;
squeal_samples[14]=40935;
squeal_samples[15]=36568;
squeal_samples[16]=32491;
squeal_samples[17]=28681;
squeal_samples[18]=25104;
squeal_samples[19]=21763;
squeal_samples[20]=18638;
squeal_samples[21]=15718;
squeal_samples[22]=12984;
squeal_samples[23]=10434;
squeal_samples[24]=8432;
squeal_samples[25]=10630;
squeal_samples[26]=13794;
squeal_samples[27]=16834;
squeal_samples[28]=19747;
squeal_samples[29]=22530;
squeal_samples[30]=25199;
squeal_samples[31]=27749;
squeal_samples[32]=30188;
squeal_samples[33]=32512;
squeal_samples[34]=34743;
squeal_samples[35]=36871;
squeal_samples[36]=38908;
squeal_samples[37]=40851;
squeal_samples[38]=42710;
squeal_samples[39]=44485;
squeal_samples[40]=46283;
squeal_samples[41]=48002;
squeal_samples[42]=49541;
squeal_samples[43]=50551;
squeal_samples[44]=46801;
squeal_samples[45]=42060;
squeal_samples[46]=37630;
squeal_samples[47]=33486;
squeal_samples[48]=29607;
squeal_samples[49]=25977;
squeal_samples[50]=22576;
squeal_samples[51]=19401;
squeal_samples[52]=16428;
squeal_samples[53]=13650;
squeal_samples[54]=11051;
squeal_samples[55]=8671;
squeal_samples[56]=9813;
squeal_samples[57]=13013;
squeal_samples[58]=16090;
squeal_samples[59]=19037;
squeal_samples[60]=21846;
squeal_samples[61]=24550;
squeal_samples[62]=27124;
squeal_samples[63]=29593;
squeal_samples[64]=31941;
squeal_samples[65]=34198;
squeal_samples[66]=36349;
squeal_samples[67]=38411;
squeal_samples[68]=40374;
squeal_samples[69]=42253;
squeal_samples[70]=44053;
squeal_samples[71]=45766;
squeal_samples[72]=47412;
squeal_samples[73]=48975;
squeal_samples[74]=50474;
squeal_samples[75]=48667;
squeal_samples[76]=43803;
squeal_samples[77]=39270;
squeal_samples[78]=35007;
squeal_samples[79]=31036;
squeal_samples[80]=27309;
squeal_samples[81]=23833;
squeal_samples[82]=20574;
squeal_samples[83]=17526;
squeal_samples[84]=14678;
squeal_samples[85]=12007;
squeal_samples[86]=9520;
squeal_samples[87]=8757;
squeal_samples[88]=11836;
squeal_samples[89]=14955;
squeal_samples[90]=17950;
squeal_samples[91]=20810;
squeal_samples[92]=23554;
squeal_samples[93]=26177;
squeal_samples[94]=28686;
squeal_samples[95]=30932;
squeal_samples[96]=33088;
squeal_samples[97]=35293;
squeal_samples[98]=37397;
squeal_samples[99]=39412;
squeal_samples[100]=41326;
squeal_samples[101]=43175;
squeal_samples[102]=44923;
squeal_samples[103]=46602;
squeal_samples[104]=48201;
squeal_samples[105]=49741;
squeal_samples[106]=50379;
squeal_samples[107]=46200;
squeal_samples[108]=41500;
squeal_samples[109]=37110;
squeal_samples[110]=32991;
squeal_samples[111]=29148;
squeal_samples[112]=25543;
squeal_samples[113]=22185;
squeal_samples[114]=19021;
squeal_samples[115]=16086;
squeal_samples[116]=13320;
squeal_samples[117]=10748;
squeal_samples[118]=8517;
squeal_samples[119]=10230;
squeal_samples[120]=13417;
squeal_samples[121]=16476;
squeal_samples[122]=19396;
squeal_samples[123]=22203;
squeal_samples[124]=24879;
squeal_samples[125]=27456;
squeal_samples[126]=29895;
squeal_samples[127]=32244;
squeal_samples[128]=34478;
squeal_samples[129]=36625;
squeal_samples[130]=38666;
squeal_samples[131]=40623;
squeal_samples[132]=42497;
squeal_samples[133]=44275;
squeal_samples[134]=45988;
squeal_samples[135]=47610;
squeal_samples[136]=49179;
squeal_samples[137]=50610;
squeal_samples[138]=48052;
squeal_samples[139]=43225;
squeal_samples[140]=38728;
squeal_samples[141]=34500;
squeal_samples[142]=30572;
squeal_samples[143]=26871;
squeal_samples[144]=23423;
squeal_samples[145]=20186;
squeal_samples[146]=17162;
squeal_samples[147]=14346;
squeal_samples[148]=11691;
squeal_samples[149]=9230;
squeal_samples[150]=9046;
squeal_samples[151]=12240;
squeal_samples[152]=15349;
squeal_samples[153]=18317;
squeal_samples[154]=21173;
squeal_samples[155]=23896;
squeal_samples[156]=26504;
squeal_samples[157]=28995;
squeal_samples[158]=31374;
squeal_samples[159]=33653;
squeal_samples[160]=35831;
squeal_samples[161]=37916;
squeal_samples[162]=39900;
squeal_samples[163]=41806;
squeal_samples[164]=43621;
squeal_samples[165]=45356;
squeal_samples[166]=47012;
squeal_samples[167]=48600;
squeal_samples[168]=50113;
squeal_samples[169]=49731;
squeal_samples[170]=45000;
squeal_samples[171]=40384;
squeal_samples[172]=36057;
squeal_samples[173]=32017;
squeal_samples[174]=28223;
squeal_samples[175]=24692;
squeal_samples[176]=21372;
squeal_samples[177]=18276;
squeal_samples[178]=15380;
squeal_samples[179]=12669;
squeal_samples[180]=10135;
squeal_samples[181]=8469;
squeal_samples[182]=11040;
squeal_samples[183]=14202;
squeal_samples[184]=17218;
squeal_samples[185]=20122;
squeal_samples[186]=22884;
squeal_samples[187]=25540;
squeal_samples[188]=28071;
squeal_samples[189]=30501;
squeal_samples[190]=32811;
squeal_samples[191]=35028;
squeal_samples[192]=37144;
squeal_samples[193]=39170;
squeal_samples[194]=41103;
squeal_samples[195]=42948;
squeal_samples[196]=44714;
squeal_samples[197]=46403;
squeal_samples[198]=48012;
squeal_samples[199]=49554;
squeal_samples[200]=50818;
squeal_samples[201]=47603;
squeal_samples[202]=42805;
squeal_samples[203]=38334;
squeal_samples[204]=34138;
squeal_samples[205]=30223;
squeal_samples[206]=26547;
squeal_samples[207]=23120;
squeal_samples[208]=19711;
squeal_samples[209]=16544;
squeal_samples[210]=13752;
squeal_samples[211]=11154;
squeal_samples[212]=8714;
squeal_samples[213]=9212;
squeal_samples[214]=12440;
squeal_samples[215]=15538;
squeal_samples[216]=18505;
squeal_samples[217]=21341;
squeal_samples[218]=24067;
squeal_samples[219]=26663;
squeal_samples[220]=29154;
squeal_samples[221]=31523;
squeal_samples[222]=33794;
squeal_samples[223]=35964;
squeal_samples[224]=38045;
squeal_samples[225]=40026;
squeal_samples[226]=41920;
squeal_samples[227]=43729;
squeal_samples[228]=45463;
squeal_samples[229]=47111;
squeal_samples[230]=48700;
squeal_samples[231]=50198;
squeal_samples[232]=49819;
squeal_samples[233]=45077;
squeal_samples[234]=40457;
squeal_samples[235]=36127;
squeal_samples[236]=32075;
squeal_samples[237]=28290;
squeal_samples[238]=24743;
squeal_samples[239]=21429;
squeal_samples[240]=18321;
squeal_samples[241]=15430;
squeal_samples[242]=12704;
squeal_samples[243]=10180;
squeal_samples[244]=8497;
squeal_samples[245]=11081;
squeal_samples[246]=14227;
squeal_samples[247]=17254;
squeal_samples[248]=20145;
squeal_samples[249]=22915;
squeal_samples[250]=25566;
squeal_samples[251]=28100;
squeal_samples[252]=30522;
squeal_samples[253]=32834;
squeal_samples[254]=35050;
squeal_samples[255]=37165;
squeal_samples[256]=39187;
squeal_samples[257]=41119;
squeal_samples[258]=42963;
squeal_samples[259]=44732;
squeal_samples[260]=46412;
squeal_samples[261]=48029;
squeal_samples[262]=49567;
squeal_samples[263]=50832;
squeal_samples[264]=47606;
squeal_samples[265]=42824;
squeal_samples[266]=38335;
squeal_samples[267]=34148;
squeal_samples[268]=30224;
squeal_samples[269]=26551;
squeal_samples[270]=23126;
squeal_samples[271]=19902;
squeal_samples[272]=16908;
squeal_samples[273]=14091;
squeal_samples[274]=11469;
squeal_samples[275]=9010;
squeal_samples[276]=8847;
squeal_samples[277]=12039;
squeal_samples[278]=15156;
squeal_samples[279]=18137;
squeal_samples[280]=20993;
squeal_samples[281]=23726;
squeal_samples[282]=26341;
squeal_samples[283]=28839;
squeal_samples[284]=31229;
squeal_samples[285]=33511;
squeal_samples[286]=35699;
squeal_samples[287]=37781;
squeal_samples[288]=39781;
squeal_samples[289]=41682;
squeal_samples[290]=43502;
squeal_samples[291]=45247;
squeal_samples[292]=46907;
squeal_samples[293]=48496;
squeal_samples[294]=50014;
squeal_samples[295]=50190;
squeal_samples[296]=45673;
squeal_samples[297]=41009;
squeal_samples[298]=36646;
squeal_samples[299]=32556;
squeal_samples[300]=28744;
squeal_samples[301]=25165;
squeal_samples[302]=21823;
squeal_samples[303]=18697;
squeal_samples[304]=15763;
squeal_samples[305]=13032;
squeal_samples[306]=10473;
squeal_samples[307]=8472;
squeal_samples[308]=10667;
squeal_samples[309]=13829;
squeal_samples[310]=16873;
squeal_samples[311]=19779;
squeal_samples[312]=22568;
squeal_samples[313]=25227;
squeal_samples[314]=27778;
squeal_samples[315]=30217;
squeal_samples[316]=32539;
squeal_samples[317]=34766;
squeal_samples[318]=36892;
squeal_samples[319]=38929;
squeal_samples[320]=40872;
squeal_samples[321]=42730;
squeal_samples[322]=44498;
squeal_samples[323]=46196;
squeal_samples[324]=47811;
squeal_samples[325]=49364;
squeal_samples[326]=50791;
squeal_samples[327]=48213;
squeal_samples[328]=43390;
squeal_samples[329]=38864;
squeal_samples[330]=34646;
squeal_samples[331]=30683;
squeal_samples[332]=26995;
squeal_samples[333]=23521;
squeal_samples[334]=20284;
squeal_samples[335]=17254;
squeal_samples[336]=14418;
squeal_samples[337]=11776;
squeal_samples[338]=9292;
squeal_samples[339]=9114;
squeal_samples[340]=12296;
squeal_samples[341]=15400;
squeal_samples[342]=18372;
squeal_samples[343]=21216;
squeal_samples[344]=23937;
squeal_samples[345]=26543;
squeal_samples[346]=29036;
squeal_samples[347]=31405;
squeal_samples[348]=33690;
squeal_samples[349]=35859;
squeal_samples[350]=37946;
squeal_samples[351]=39928;
squeal_samples[352]=41823;
squeal_samples[353]=43640;
squeal_samples[354]=45367;
squeal_samples[355]=47029;
squeal_samples[356]=48607;
squeal_samples[357]=50122;
squeal_samples[358]=50292;
squeal_samples[359]=45769;
squeal_samples[360]=41097;
squeal_samples[361]=36722;
squeal_samples[362]=32634;
squeal_samples[363]=28811;
squeal_samples[364]=25229;
squeal_samples[365]=21882;
squeal_samples[366]=18746;
squeal_samples[367]=15813;
squeal_samples[368]=13078;
squeal_samples[369]=10508;
squeal_samples[370]=8509;
squeal_samples[371]=10695;
squeal_samples[372]=13861;
squeal_samples[373]=16902;
squeal_samples[374]=19803;
squeal_samples[375]=22593;
squeal_samples[376]=25250;
squeal_samples[377]=27800;
squeal_samples[378]=30231;
squeal_samples[379]=32562;
squeal_samples[380]=34774;
squeal_samples[381]=36909;
squeal_samples[382]=38940;
squeal_samples[383]=40880;
squeal_samples[384]=42736;
squeal_samples[385]=44506;
squeal_samples[386]=46201;
squeal_samples[387]=47820;
squeal_samples[388]=49365;
squeal_samples[389]=50795;
squeal_samples[390]=48217;
squeal_samples[391]=43387;
squeal_samples[392]=38870;
squeal_samples[393]=34636;
squeal_samples[394]=30683;
squeal_samples[395]=26980;
squeal_samples[396]=23514;
squeal_samples[397]=20277;
squeal_samples[398]=17249;
squeal_samples[399]=14409;
squeal_samples[400]=11762;
squeal_samples[401]=9284;
squeal_samples[402]=9095;
squeal_samples[403]=12287;
squeal_samples[404]=15387;
squeal_samples[405]=18362;
squeal_samples[406]=21196;
squeal_samples[407]=23930;
squeal_samples[408]=26523;
squeal_samples[409]=29019;
squeal_samples[410]=31395;
squeal_samples[411]=33668;
squeal_samples[412]=35848;
squeal_samples[413]=37923;
squeal_samples[414]=39913;
squeal_samples[415]=41805;
squeal_samples[416]=43621;
squeal_samples[417]=45350;
squeal_samples[418]=47010;
squeal_samples[419]=48589;
squeal_samples[420]=50104;
squeal_samples[421]=50274;
squeal_samples[422]=45749;
squeal_samples[423]=41079;
squeal_samples[424]=36704;
squeal_samples[425]=32614;
squeal_samples[426]=28792;
squeal_samples[427]=25206;
squeal_samples[428]=21855;
squeal_samples[429]=18725;
squeal_samples[430]=15786;
squeal_samples[431]=13053;
squeal_samples[432]=10489;
squeal_samples[433]=8490;
squeal_samples[434]=10673;
squeal_samples[435]=13840;
squeal_samples[436]=16872;
squeal_samples[437]=19782;
squeal_samples[438]=22563;
squeal_samples[439]=25229;
squeal_samples[440]=27769;
squeal_samples[441]=30211;
squeal_samples[442]=32530;
squeal_samples[443]=34759;
squeal_samples[444]=36878;
squeal_samples[445]=38918;
squeal_samples[446]=40850;
squeal_samples[447]=42712;
squeal_samples[448]=44483;
squeal_samples[449]=46177;
squeal_samples[450]=47790;
squeal_samples[451]=49346;
squeal_samples[452]=50768;
squeal_samples[453]=48189;
squeal_samples[454]=43362;
squeal_samples[455]=38840;
squeal_samples[456]=34610;
squeal_samples[457]=30656;
squeal_samples[458]=26953;
squeal_samples[459]=23490;
squeal_samples[460]=20253;
squeal_samples[461]=17216;
squeal_samples[462]=14385;
squeal_samples[463]=11733;
squeal_samples[464]=9255;
squeal_samples[465]=9069;
squeal_samples[466]=12256;
squeal_samples[467]=15361;
squeal_samples[468]=18331;
squeal_samples[469]=21172;
squeal_samples[470]=23897;
squeal_samples[471]=26497;
squeal_samples[472]=28989;
squeal_samples[473]=31366;
squeal_samples[474]=33640;
squeal_samples[475]=35818;
squeal_samples[476]=37895;
squeal_samples[477]=39883;
squeal_samples[478]=41776;
squeal_samples[479]=43591;
squeal_samples[480]=45322;
squeal_samples[481]=46979;
squeal_samples[482]=48561;
squeal_samples[483]=50072;
squeal_samples[484]=50245;
squeal_samples[485]=45721;
squeal_samples[486]=41047;
squeal_samples[487]=36675;
squeal_samples[488]=32583;
squeal_samples[489]=28763;
squeal_samples[490]=25174;
squeal_samples[491]=21827;
squeal_samples[492]=18691;
squeal_samples[493]=15758;
squeal_samples[494]=13021;
squeal_samples[495]=10460;
squeal_samples[496]=8456;
squeal_samples[497]=10647;
squeal_samples[498]=13802;
squeal_samples[499]=16848;
squeal_samples[500]=19744;
squeal_samples[501]=22539;
squeal_samples[502]=25191;
squeal_samples[503]=27742;
squeal_samples[504]=30177;
squeal_samples[505]=32499;
squeal_samples[506]=34728;
squeal_samples[507]=36846;
squeal_samples[508]=38884;
squeal_samples[509]=40822;
squeal_samples[510]=42676;
squeal_samples[511]=44454;
squeal_samples[512]=46142;
squeal_samples[513]=47760;
squeal_samples[514]=49312;
squeal_samples[515]=50737;
squeal_samples[516]=48156;
squeal_samples[517]=43328;
squeal_samples[518]=38810;
squeal_samples[519]=34575;
squeal_samples[520]=30624;
squeal_samples[521]=26919;
squeal_samples[522]=23458;
squeal_samples[523]=20219;
squeal_samples[524]=17184;
squeal_samples[525]=14351;
squeal_samples[526]=11699;
squeal_samples[527]=9223;
squeal_samples[528]=9034;
squeal_samples[529]=12223;
squeal_samples[530]=15328;
squeal_samples[531]=18296;
squeal_samples[532]=21139;
squeal_samples[533]=23862;
squeal_samples[534]=26464;
squeal_samples[535]=28955;
squeal_samples[536]=31331;
squeal_samples[537]=33607;
squeal_samples[538]=35782;
squeal_samples[539]=37863;
squeal_samples[540]=39846;
squeal_samples[541]=41744;
squeal_samples[542]=43554;
squeal_samples[543]=45289;
squeal_samples[544]=46943;
squeal_samples[545]=48527;
squeal_samples[546]=50038;
squeal_samples[547]=50208;
squeal_samples[548]=45688;
squeal_samples[549]=41009;
squeal_samples[550]=36643;
squeal_samples[551]=32545;
squeal_samples[552]=28730;
squeal_samples[553]=25136;
squeal_samples[554]=21794;
squeal_samples[555]=18653;
squeal_samples[556]=15725;
squeal_samples[557]=12983;
squeal_samples[558]=10425;
squeal_samples[559]=8421;
squeal_samples[560]=10608;
squeal_samples[561]=13770;
squeal_samples[562]=16808;
squeal_samples[563]=19712;
squeal_samples[564]=22499;
squeal_samples[565]=25156;
squeal_samples[566]=27706;
squeal_samples[567]=30138;
squeal_samples[568]=32466;
squeal_samples[569]=34688;
squeal_samples[570]=36812;
squeal_samples[571]=38845;
squeal_samples[572]=40786;
squeal_samples[573]=42638;
squeal_samples[574]=44419;
squeal_samples[575]=46102;
squeal_samples[576]=47725;
squeal_samples[577]=49272;
squeal_samples[578]=50749;
squeal_samples[579]=48918;
squeal_samples[580]=44034;
squeal_samples[581]=39468;
squeal_samples[582]=35189;
squeal_samples[583]=31196;
squeal_samples[584]=27454;
squeal_samples[585]=23957;
squeal_samples[586]=20675;
squeal_samples[587]=17620;
squeal_samples[588]=14743;
squeal_samples[589]=12077;
squeal_samples[590]=9565;
squeal_samples[591]=8317;
squeal_samples[592]=11191;
squeal_samples[593]=14332;
squeal_samples[594]=17342;
squeal_samples[595]=20226;
squeal_samples[596]=22987;
squeal_samples[597]=25628;
squeal_samples[598]=28149;
squeal_samples[599]=30567;
squeal_samples[600]=32867;
squeal_samples[601]=35078;
squeal_samples[602]=37178;
squeal_samples[603]=39200;
squeal_samples[604]=41118;
squeal_samples[605]=42966;
squeal_samples[606]=44714;
squeal_samples[607]=46395;
squeal_samples[608]=48003;
squeal_samples[609]=49535;
squeal_samples[610]=50795;
squeal_samples[611]=47564;
squeal_samples[612]=42766;
squeal_samples[613]=38279;
squeal_samples[614]=34077;
squeal_samples[615]=30160;
squeal_samples[616]=26477;
squeal_samples[617]=23041;
squeal_samples[618]=19818;
squeal_samples[619]=16815;
squeal_samples[620]=13997;
squeal_samples[621]=11368;
squeal_samples[622]=8905;
squeal_samples[623]=9380;
squeal_samples[624]=12597;
squeal_samples[625]=15678;
squeal_samples[626]=18636;
squeal_samples[627]=21458;
squeal_samples[628]=24167;
squeal_samples[629]=26753;
squeal_samples[630]=29225;
squeal_samples[631]=31587;
squeal_samples[632]=33851;
squeal_samples[633]=36009;
squeal_samples[634]=38081;
squeal_samples[635]=40046;
squeal_samples[636]=41939;
squeal_samples[637]=43738;
squeal_samples[638]=45461;
squeal_samples[639]=47107;
squeal_samples[640]=48677;
squeal_samples[641]=50177;
squeal_samples[642]=50340;
squeal_samples[643]=45802;
squeal_samples[644]=41122;
squeal_samples[645]=36734;
squeal_samples[646]=32635;
squeal_samples[647]=28799;
squeal_samples[648]=25211;
squeal_samples[649]=21848;
squeal_samples[650]=18708;
squeal_samples[651]=15771;
squeal_samples[652]=13019;
squeal_samples[653]=10455;
squeal_samples[654]=8448;
squeal_samples[655]=10626;
squeal_samples[656]=13791;
squeal_samples[657]=16822;
squeal_samples[658]=19725;
squeal_samples[659]=22507;
squeal_samples[660]=25161;
squeal_samples[661]=27707;
squeal_samples[662]=30137;
squeal_samples[663]=32458;
squeal_samples[664]=34679;
squeal_samples[665]=36803;
squeal_samples[666]=38834;
squeal_samples[667]=40769;
squeal_samples[668]=42627;
squeal_samples[669]=44397;
squeal_samples[670]=46084;
squeal_samples[671]=47705;
squeal_samples[672]=49248;
squeal_samples[673]=50723;
squeal_samples[674]=48887;
squeal_samples[675]=44004;
squeal_samples[676]=39436;
squeal_samples[677]=35161;
squeal_samples[678]=31156;
squeal_samples[679]=27415;
squeal_samples[680]=23912;
squeal_samples[681]=20635;
squeal_samples[682]=17577;
squeal_samples[683]=14700;
squeal_samples[684]=12030;
squeal_samples[685]=9515;
squeal_samples[686]=8749;
squeal_samples[687]=11809;
squeal_samples[688]=14928;
squeal_samples[689]=17910;
squeal_samples[690]=20771;
squeal_samples[691]=23497;
squeal_samples[692]=26119;
squeal_samples[693]=28615;
squeal_samples[694]=31004;
squeal_samples[695]=33283;
squeal_samples[696]=35474;
squeal_samples[697]=37557;
squeal_samples[698]=39553;
squeal_samples[699]=41461;
squeal_samples[700]=43275;
squeal_samples[701]=45023;
squeal_samples[702]=46680;
squeal_samples[703]=48271;
squeal_samples[704]=49789;
squeal_samples[705]=50780;
squeal_samples[706]=46997;
squeal_samples[707]=42240;
squeal_samples[708]=37778;
squeal_samples[709]=33605;
squeal_samples[710]=29708;
squeal_samples[711]=26054;
squeal_samples[712]=22642;
squeal_samples[713]=19440;
squeal_samples[714]=16454;
squeal_samples[715]=13655;
squeal_samples[716]=11047;
squeal_samples[717]=8646;
squeal_samples[718]=9781;
squeal_samples[719]=12970;
squeal_samples[720]=16042;
squeal_samples[721]=18973;
squeal_samples[722]=21785;
squeal_samples[723]=24470;
squeal_samples[724]=27043;
squeal_samples[725]=29501;
squeal_samples[726]=31849;
squeal_samples[727]=34091;
squeal_samples[728]=36244;
squeal_samples[729]=38294;
squeal_samples[730]=40257;
squeal_samples[731]=42134;
squeal_samples[732]=43915;
squeal_samples[733]=45628;
squeal_samples[734]=47263;
squeal_samples[735]=48828;
squeal_samples[736]=50317;
squeal_samples[737]=49915;
squeal_samples[738]=45152;
squeal_samples[739]=40514;
squeal_samples[740]=36154;
squeal_samples[741]=32092;
squeal_samples[742]=28286;
squeal_samples[743]=24726;
squeal_samples[744]=21395;
squeal_samples[745]=18276;
squeal_samples[746]=15362;
squeal_samples[747]=12632;
squeal_samples[748]=10088;
squeal_samples[749]=8408;
squeal_samples[750]=10971;
squeal_samples[751]=14121;
squeal_samples[752]=17133;
squeal_samples[753]=20023;
squeal_samples[754]=22787;
squeal_samples[755]=25429;
squeal_samples[756]=27961;
squeal_samples[757]=30372;
squeal_samples[758]=32683;
squeal_samples[759]=34889;
squeal_samples[760]=37002;
squeal_samples[761]=39018;
squeal_samples[762]=40950;
squeal_samples[763]=42782;
squeal_samples[764]=44550;
squeal_samples[765]=46227;
squeal_samples[766]=47837;
squeal_samples[767]=49372;
squeal_samples[768]=50783;
squeal_samples[769]=48201;
squeal_samples[770]=43354;
squeal_samples[771]=38820;
squeal_samples[772]=34579;
squeal_samples[773]=30614;
squeal_samples[774]=26898;
squeal_samples[775]=23427;
squeal_samples[776]=20177;
squeal_samples[777]=17134;
squeal_samples[778]=14296;
squeal_samples[779]=11635;
squeal_samples[780]=9152;
squeal_samples[781]=8959;
squeal_samples[782]=12147;
squeal_samples[783]=15240;
squeal_samples[784]=18211;
squeal_samples[785]=21044;
squeal_samples[786]=23770;
squeal_samples[787]=26366;
squeal_samples[788]=28854;
squeal_samples[789]=31225;
squeal_samples[790]=33499;
squeal_samples[791]=35670;
squeal_samples[792]=37743;
squeal_samples[793]=39729;
squeal_samples[794]=41624;
squeal_samples[795]=43436;
squeal_samples[796]=45164;
squeal_samples[797]=46814;
squeal_samples[798]=48395;
squeal_samples[799]=49907;
squeal_samples[800]=50531;
squeal_samples[801]=46319;
squeal_samples[802]=41597;
squeal_samples[803]=37172;
squeal_samples[804]=33041;
squeal_samples[805]=29167;
squeal_samples[806]=25548;
squeal_samples[807]=22160;
squeal_samples[808]=18988;
squeal_samples[809]=16030;
squeal_samples[810]=13250;
squeal_samples[811]=10665;
squeal_samples[812]=8413;
squeal_samples[813]=10117;
squeal_samples[814]=13296;
squeal_samples[815]=16343;
squeal_samples[816]=19266;
squeal_samples[817]=22054;
squeal_samples[818]=24734;
squeal_samples[819]=27286;
squeal_samples[820]=29739;
squeal_samples[821]=32063;
squeal_samples[822]=34302;
squeal_samples[823]=36431;
squeal_samples[824]=38478;
squeal_samples[825]=40423;
squeal_samples[826]=42294;
squeal_samples[827]=44067;
squeal_samples[828]=45772;
squeal_samples[829]=47393;
squeal_samples[830]=48948;
squeal_samples[831]=50434;
squeal_samples[832]=49359;
squeal_samples[833]=44488;
squeal_samples[834]=39880;
squeal_samples[835]=35568;
squeal_samples[836]=31529;
squeal_samples[837]=27764;
squeal_samples[838]=24222;
squeal_samples[839]=20927;
squeal_samples[840]=17830;
squeal_samples[841]=14940;
squeal_samples[842]=12235;
squeal_samples[843]=9709;
squeal_samples[844]=8440;
squeal_samples[845]=11299;
squeal_samples[846]=14432;
squeal_samples[847]=17425;
squeal_samples[848]=20303;
squeal_samples[849]=23051;
squeal_samples[850]=25681;
squeal_samples[851]=28194;
squeal_samples[852]=30591;
squeal_samples[853]=32894;
squeal_samples[854]=35091;
squeal_samples[855]=37186;
squeal_samples[856]=39195;
squeal_samples[857]=41108;
squeal_samples[858]=42946;
squeal_samples[859]=44693;
squeal_samples[860]=46365;
squeal_samples[861]=47964;
squeal_samples[862]=49488;
squeal_samples[863]=50745;
squeal_samples[864]=47502;
squeal_samples[865]=42700;
squeal_samples[866]=38205;
squeal_samples[867]=34000;
squeal_samples[868]=30068;
squeal_samples[869]=26386;
squeal_samples[870]=22937;
squeal_samples[871]=19717;
squeal_samples[872]=16699;
squeal_samples[873]=13884;
squeal_samples[874]=11243;
squeal_samples[875]=8785;
squeal_samples[876]=9251;
squeal_samples[877]=12469;
squeal_samples[878]=15546;
squeal_samples[879]=18501;
squeal_samples[880]=21326;
squeal_samples[881]=24027;
squeal_samples[882]=26614;
squeal_samples[883]=29086;
squeal_samples[884]=31443;
squeal_samples[885]=33705;
squeal_samples[886]=35867;
squeal_samples[887]=37927;
squeal_samples[888]=39898;
squeal_samples[889]=41782;
squeal_samples[890]=43583;
squeal_samples[891]=45306;
squeal_samples[892]=46949;
squeal_samples[893]=48523;
squeal_samples[894]=50019;
squeal_samples[895]=50181;
squeal_samples[896]=45639;
squeal_samples[897]=40961;
squeal_samples[898]=36572;
squeal_samples[899]=32468;
squeal_samples[900]=28632;
squeal_samples[901]=25044;
squeal_samples[902]=21680;
squeal_samples[903]=18535;
squeal_samples[904]=15598;
squeal_samples[905]=12846;
squeal_samples[906]=10284;
squeal_samples[907]=8272;
squeal_samples[908]=10455;
squeal_samples[909]=13617;
squeal_samples[910]=16648;
squeal_samples[911]=19548;
squeal_samples[912]=22327;
squeal_samples[913]=24989;
squeal_samples[914]=27527;
squeal_samples[915]=29961;
squeal_samples[916]=32280;
squeal_samples[917]=34504;
squeal_samples[918]=36623;
squeal_samples[919]=38654;
squeal_samples[920]=40591;
squeal_samples[921]=42448;
squeal_samples[922]=44217;
squeal_samples[923]=45907;
squeal_samples[924]=47518;
squeal_samples[925]=49070;
squeal_samples[926]=50543;
squeal_samples[927]=48708;
squeal_samples[928]=43826;
squeal_samples[929]=39254;
squeal_samples[930]=34979;
squeal_samples[931]=30974;
squeal_samples[932]=27239;
squeal_samples[933]=23730;
squeal_samples[934]=20452;
squeal_samples[935]=17389;
squeal_samples[936]=14519;
squeal_samples[937]=11842;
squeal_samples[938]=9333;
squeal_samples[939]=8561;
squeal_samples[940]=11632;
squeal_samples[941]=14746;
squeal_samples[942]=17727;
squeal_samples[943]=20584;
squeal_samples[944]=23315;
squeal_samples[945]=25930;
squeal_samples[946]=28433;
squeal_samples[947]=30815;
squeal_samples[948]=33101;
squeal_samples[949]=35289;
squeal_samples[950]=37375;
squeal_samples[951]=39371;
squeal_samples[952]=41271;
squeal_samples[953]=43099;
squeal_samples[954]=44835;
squeal_samples[955]=46496;
squeal_samples[956]=48090;
squeal_samples[957]=49603;
squeal_samples[958]=50855;
squeal_samples[959]=47600;
squeal_samples[960]=42788;
squeal_samples[961]=38280;
squeal_samples[962]=34070;
squeal_samples[963]=30119;
squeal_samples[964]=26441;
squeal_samples[965]=22976;
squeal_samples[966]=19755;
squeal_samples[967]=16726;
squeal_samples[968]=13907;
squeal_samples[969]=11262;
squeal_samples[970]=8794;
squeal_samples[971]=9261;
squeal_samples[972]=12473;
squeal_samples[973]=15550;
squeal_samples[974]=18496;
squeal_samples[975]=21323;
squeal_samples[976]=24016;
squeal_samples[977]=26606;
squeal_samples[978]=29069;
squeal_samples[979]=31431;
squeal_samples[980]=33684;
squeal_samples[981]=35846;
squeal_samples[982]=37908;
squeal_samples[983]=39878;
squeal_samples[984]=41755;
squeal_samples[985]=43561;
squeal_samples[986]=45270;
squeal_samples[987]=46918;
squeal_samples[988]=48482;
squeal_samples[989]=49987;
squeal_samples[990]=50142;
squeal_samples[991]=45599;
squeal_samples[992]=40918;
squeal_samples[993]=36526;
squeal_samples[994]=32427;
squeal_samples[995]=28590;
squeal_samples[996]=24997;
squeal_samples[997]=21632;
squeal_samples[998]=18492;
squeal_samples[999]=15542;
squeal_samples[1000]=12798;
squeal_samples[1001]=10223;
squeal_samples[1002]=8216;
squeal_samples[1003]=10397;
squeal_samples[1004]=13561;
squeal_samples[1005]=16588;
squeal_samples[1006]=19500;
squeal_samples[1007]=22267;
squeal_samples[1008]=24932;
squeal_samples[1009]=27471;
squeal_samples[1010]=29901;
squeal_samples[1011]=32227;
squeal_samples[1012]=34443;
squeal_samples[1013]=36567;
squeal_samples[1014]=38598;
squeal_samples[1015]=40532;
squeal_samples[1016]=42388;
squeal_samples[1017]=44151;
squeal_samples[1018]=45847;
squeal_samples[1019]=47460;
squeal_samples[1020]=49007;
squeal_samples[1021]=50481;
squeal_samples[1022]=49399;
squeal_samples[1023]=44515;
squeal_samples[1024]=39893;
squeal_samples[1025]=35578;
squeal_samples[1026]=31527;
squeal_samples[1027]=27751;
squeal_samples[1028]=24205;
squeal_samples[1029]=20897;
squeal_samples[1030]=17798;
squeal_samples[1031]=14898;
squeal_samples[1032]=12192;
squeal_samples[1033]=9658;
squeal_samples[1034]=8385;
squeal_samples[1035]=11237;
squeal_samples[1036]=14372;
squeal_samples[1037]=17357;
squeal_samples[1038]=20239;
squeal_samples[1039]=22972;
squeal_samples[1040]=25607;
squeal_samples[1041]=28113;
squeal_samples[1042]=30518;
squeal_samples[1043]=32808;
squeal_samples[1044]=35007;
squeal_samples[1045]=37095;
squeal_samples[1046]=39111;
squeal_samples[1047]=41012;
squeal_samples[1048]=42851;
squeal_samples[1049]=44591;
squeal_samples[1050]=46269;
squeal_samples[1051]=47864;
squeal_samples[1052]=49386;
squeal_samples[1053]=50797;
squeal_samples[1054]=48193;
squeal_samples[1055]=43335;
squeal_samples[1056]=38791;
squeal_samples[1057]=34539;
squeal_samples[1058]=30556;
squeal_samples[1059]=26842;
squeal_samples[1060]=23356;
squeal_samples[1061]=20096;
squeal_samples[1062]=17050;
squeal_samples[1063]=14197;
squeal_samples[1064]=11533;
squeal_samples[1065]=9045;
squeal_samples[1066]=8840;
squeal_samples[1067]=12029;
squeal_samples[1068]=15117;
squeal_samples[1069]=18086;
squeal_samples[1070]=20917;
squeal_samples[1071]=23633;
squeal_samples[1072]=26235;
squeal_samples[1073]=28710;
squeal_samples[1074]=31091;
squeal_samples[1075]=33349;
squeal_samples[1076]=35529;
squeal_samples[1077]=37595;
squeal_samples[1078]=39581;
squeal_samples[1079]=41467;
squeal_samples[1080]=43276;
squeal_samples[1081]=45008;
squeal_samples[1082]=46659;
squeal_samples[1083]=48234;
squeal_samples[1084]=49740;
squeal_samples[1085]=50723;
squeal_samples[1086]=46932;
squeal_samples[1087]=42157;
squeal_samples[1088]=37683;
squeal_samples[1089]=33502;
squeal_samples[1090]=29590;
squeal_samples[1091]=25932;
squeal_samples[1092]=22502;
squeal_samples[1093]=19300;
squeal_samples[1094]=16299;
squeal_samples[1095]=13498;
squeal_samples[1096]=10876;
squeal_samples[1097]=8476;
squeal_samples[1098]=9594;
squeal_samples[1099]=12798;
squeal_samples[1100]=15849;
squeal_samples[1101]=18789;
squeal_samples[1102]=21591;
squeal_samples[1103]=24276;
squeal_samples[1104]=26840;
squeal_samples[1105]=29302;
squeal_samples[1106]=31639;
squeal_samples[1107]=33888;
squeal_samples[1108]=36032;
squeal_samples[1109]=38079;
squeal_samples[1110]=40045;
squeal_samples[1111]=41906;
squeal_samples[1112]=43701;
squeal_samples[1113]=45406;
squeal_samples[1114]=47038;
squeal_samples[1115]=48602;
squeal_samples[1116]=50089;
squeal_samples[1117]=50241;
squeal_samples[1118]=45687;
squeal_samples[1119]=40990;
squeal_samples[1120]=36593;
squeal_samples[1121]=32476;
squeal_samples[1122]=28633;
squeal_samples[1123]=25026;
squeal_samples[1124]=21667;
squeal_samples[1125]=18504;
squeal_samples[1126]=15565;
squeal_samples[1127]=12803;
squeal_samples[1128]=10223;
squeal_samples[1129]=8218;
squeal_samples[1130]=10388;
squeal_samples[1131]=13557;
squeal_samples[1132]=16572;
squeal_samples[1133]=19480;
squeal_samples[1134]=22248;
squeal_samples[1135]=24914;
squeal_samples[1136]=27443;
squeal_samples[1137]=29881;
squeal_samples[1138]=32193;
squeal_samples[1139]=34412;
squeal_samples[1140]=36529;
squeal_samples[1141]=38563;
squeal_samples[1142]=40493;
squeal_samples[1143]=42345;
squeal_samples[1144]=44115;
squeal_samples[1145]=45803;
squeal_samples[1146]=47416;
squeal_samples[1147]=48957;
squeal_samples[1148]=50428;
squeal_samples[1149]=49351;
squeal_samples[1150]=44462;
squeal_samples[1151]=39844;
squeal_samples[1152]=35520;
squeal_samples[1153]=31474;
squeal_samples[1154]=27687;
squeal_samples[1155]=24147;
squeal_samples[1156]=20833;
squeal_samples[1157]=17734;
squeal_samples[1158]=14835;
squeal_samples[1159]=12128;
squeal_samples[1160]=9589;
squeal_samples[1161]=8315;
squeal_samples[1162]=11172;
squeal_samples[1163]=14298;
squeal_samples[1164]=17295;
squeal_samples[1165]=20163;
squeal_samples[1166]=22911;
squeal_samples[1167]=25531;
squeal_samples[1168]=28047;
squeal_samples[1169]=30442;
squeal_samples[1170]=32742;
squeal_samples[1171]=34933;
squeal_samples[1172]=37027;
squeal_samples[1173]=39031;
squeal_samples[1174]=40946;
squeal_samples[1175]=42776;
squeal_samples[1176]=44525;
squeal_samples[1177]=46191;
squeal_samples[1178]=47788;
squeal_samples[1179]=49311;
squeal_samples[1180]=50722;
squeal_samples[1181]=48118;
squeal_samples[1182]=43258;
squeal_samples[1183]=38718;
squeal_samples[1184]=34461;
squeal_samples[1185]=30484;
squeal_samples[1186]=26760;
squeal_samples[1187]=23281;
squeal_samples[1188]=20021;
squeal_samples[1189]=16976;
squeal_samples[1190]=14121;
squeal_samples[1191]=11455;
squeal_samples[1192]=8963;
squeal_samples[1193]=8766;
squeal_samples[1194]=11949;
squeal_samples[1195]=15038;
squeal_samples[1196]=18005;
squeal_samples[1197]=20845;
squeal_samples[1198]=23557;
squeal_samples[1199]=26156;
squeal_samples[1200]=28638;
squeal_samples[1201]=31008;
squeal_samples[1202]=33273;
squeal_samples[1203]=35448;
squeal_samples[1204]=37518;
squeal_samples[1205]=39500;
squeal_samples[1206]=41396;
squeal_samples[1207]=43201;
squeal_samples[1208]=44930;
squeal_samples[1209]=46579;
squeal_samples[1210]=48157;
squeal_samples[1211]=49660;
squeal_samples[1212]=50647;
squeal_samples[1213]=46852;
squeal_samples[1214]=42078;
squeal_samples[1215]=37606;
squeal_samples[1216]=33423;
squeal_samples[1217]=29513;
squeal_samples[1218]=25853;
squeal_samples[1219]=22425;
squeal_samples[1220]=19221;
squeal_samples[1221]=16223;
squeal_samples[1222]=13419;
squeal_samples[1223]=10801;
squeal_samples[1224]=8394;
squeal_samples[1225]=9522;
squeal_samples[1226]=12717;
squeal_samples[1227]=15775;
squeal_samples[1228]=18709;
squeal_samples[1229]=21516;
squeal_samples[1230]=24197;
squeal_samples[1231]=26766;
squeal_samples[1232]=29223;
squeal_samples[1233]=31564;
squeal_samples[1234]=33810;
squeal_samples[1235]=35955;
squeal_samples[1236]=38005;
squeal_samples[1237]=39966;
squeal_samples[1238]=41832;
squeal_samples[1239]=43624;
squeal_samples[1240]=45329;
squeal_samples[1241]=46965;
squeal_samples[1242]=48522;
squeal_samples[1243]=50017;
squeal_samples[1244]=50162;
squeal_samples[1245]=45615;
squeal_samples[1246]=40911;
squeal_samples[1247]=36520;
squeal_samples[1248]=32399;
squeal_samples[1249]=28557;
squeal_samples[1250]=24954;
squeal_samples[1251]=21587;
squeal_samples[1252]=18434;
squeal_samples[1253]=15485;
squeal_samples[1254]=12730;
squeal_samples[1255]=10151;
squeal_samples[1256]=8137;
squeal_samples[1257]=10320;
squeal_samples[1258]=13476;
squeal_samples[1259]=16502;
squeal_samples[1260]=19402;
squeal_samples[1261]=22178;
squeal_samples[1262]=24835;
squeal_samples[1263]=27373;
squeal_samples[1264]=29804;
squeal_samples[1265]=32119;
squeal_samples[1266]=34338;
squeal_samples[1267]=36458;
squeal_samples[1268]=38486;
squeal_samples[1269]=40422;
squeal_samples[1270]=42268;
squeal_samples[1271]=44044;
squeal_samples[1272]=45729;
squeal_samples[1273]=47344;
squeal_samples[1274]=48880;
squeal_samples[1275]=50359;
squeal_samples[1276]=49274;
squeal_samples[1277]=44393;
squeal_samples[1278]=39768;
squeal_samples[1279]=35449;
squeal_samples[1280]=31398;
squeal_samples[1281]=27618;
squeal_samples[1282]=24072;
squeal_samples[1283]=20762;
squeal_samples[1284]=17660;
squeal_samples[1285]=14763;
squeal_samples[1286]=12056;
squeal_samples[1287]=9516;
squeal_samples[1288]=8245;
squeal_samples[1289]=11096;
squeal_samples[1290]=14230;
squeal_samples[1291]=17221;
squeal_samples[1292]=20092;
squeal_samples[1293]=22839;
squeal_samples[1294]=25459;
squeal_samples[1295]=27975;
squeal_samples[1296]=30372;
squeal_samples[1297]=32669;
squeal_samples[1298]=34862;
squeal_samples[1299]=36956;
squeal_samples[1300]=38960;
squeal_samples[1301]=40874;
squeal_samples[1302]=42707;
squeal_samples[1303]=44451;
squeal_samples[1304]=46123;
squeal_samples[1305]=47715;
squeal_samples[1306]=49243;
squeal_samples[1307]=50650;
squeal_samples[1308]=48046;
squeal_samples[1309]=43191;
squeal_samples[1310]=38643;
squeal_samples[1311]=34396;
squeal_samples[1312]=30409;
squeal_samples[1313]=26694;
squeal_samples[1314]=23208;
squeal_samples[1315]=19953;
squeal_samples[1316]=16904;
squeal_samples[1317]=14053;
squeal_samples[1318]=11385;
squeal_samples[1319]=8893;
squeal_samples[1320]=8698;
squeal_samples[1321]=11878;
squeal_samples[1322]=14969;
squeal_samples[1323]=17936;
squeal_samples[1324]=20773;
squeal_samples[1325]=23493;
squeal_samples[1326]=26083;
squeal_samples[1327]=28571;
squeal_samples[1328]=30937;
squeal_samples[1329]=33205;
squeal_samples[1330]=35380;
squeal_samples[1331]=37448;
squeal_samples[1332]=39433;
squeal_samples[1333]=41325;
squeal_samples[1334]=43133;
squeal_samples[1335]=44863;
squeal_samples[1336]=46509;
squeal_samples[1337]=48089;
squeal_samples[1338]=49592;
squeal_samples[1339]=50832;
squeal_samples[1340]=47567;
squeal_samples[1341]=42745;
squeal_samples[1342]=38226;
squeal_samples[1343]=34002;
squeal_samples[1344]=30050;
squeal_samples[1345]=26346;
squeal_samples[1346]=22888;
squeal_samples[1347]=19645;
squeal_samples[1348]=16618;
squeal_samples[1349]=13782;
squeal_samples[1350]=11133;
squeal_samples[1351]=8662;
squeal_samples[1352]=9119;
squeal_samples[1353]=12332;
squeal_samples[1354]=15403;
squeal_samples[1355]=18349;
squeal_samples[1356]=21166;
squeal_samples[1357]=23865;
squeal_samples[1358]=26443;
squeal_samples[1359]=28914;
squeal_samples[1360]=31263;
squeal_samples[1361]=33522;
squeal_samples[1362]=35675;
squeal_samples[1363]=37735;
squeal_samples[1364]=39701;
squeal_samples[1365]=41585;
squeal_samples[1366]=43376;
squeal_samples[1367]=45096;
squeal_samples[1368]=46735;
squeal_samples[1369]=48299;
squeal_samples[1370]=49797;
squeal_samples[1371]=50765;
squeal_samples[1372]=46967;
squeal_samples[1373]=42173;
squeal_samples[1374]=37690;
squeal_samples[1375]=33499;
squeal_samples[1376]=29580;
squeal_samples[1377]=25912;
squeal_samples[1378]=22472;
squeal_samples[1379]=19258;
squeal_samples[1380]=16254;
squeal_samples[1381]=13446;
squeal_samples[1382]=10812;
squeal_samples[1383]=8410;
squeal_samples[1384]=9525;
squeal_samples[1385]=12723;
squeal_samples[1386]=15768;
squeal_samples[1387]=18709;
squeal_samples[1388]=21498;
squeal_samples[1389]=24191;
squeal_samples[1390]=26752;
squeal_samples[1391]=29207;
squeal_samples[1392]=31549;
squeal_samples[1393]=33786;
squeal_samples[1394]=35935;
squeal_samples[1395]=37978;
squeal_samples[1396]=39933;
squeal_samples[1397]=41805;
squeal_samples[1398]=43587;
squeal_samples[1399]=45297;
squeal_samples[1400]=46926;
squeal_samples[1401]=48481;
squeal_samples[1402]=49971;
squeal_samples[1403]=50579;
squeal_samples[1404]=46335;
squeal_samples[1405]=41590;
squeal_samples[1406]=37141;
squeal_samples[1407]=32986;
squeal_samples[1408]=29098;
squeal_samples[1409]=25457;
squeal_samples[1410]=22050;
squeal_samples[1411]=18863;
squeal_samples[1412]=15882;
squeal_samples[1413]=13091;
squeal_samples[1414]=10494;
squeal_samples[1415]=8224;
squeal_samples[1416]=9927;
squeal_samples[1417]=13090;
squeal_samples[1418]=16138;
squeal_samples[1419]=19044;
squeal_samples[1420]=21839;
squeal_samples[1421]=24502;
squeal_samples[1422]=27054;
squeal_samples[1423]=29493;
squeal_samples[1424]=31818;
squeal_samples[1425]=34055;
squeal_samples[1426]=36173;
squeal_samples[1427]=38220;
squeal_samples[1428]=40152;
squeal_samples[1429]=42023;
squeal_samples[1430]=43793;
squeal_samples[1431]=45490;
squeal_samples[1432]=47112;
squeal_samples[1433]=48659;
squeal_samples[1434]=50139;
squeal_samples[1435]=50278;
squeal_samples[1436]=45714;
squeal_samples[1437]=41001;
squeal_samples[1438]=36600;
squeal_samples[1439]=32466;
squeal_samples[1440]=28616;
squeal_samples[1441]=25001;
squeal_samples[1442]=21623;
squeal_samples[1443]=18464;
squeal_samples[1444]=15507;
squeal_samples[1445]=12745;
squeal_samples[1446]=10159;
squeal_samples[1447]=8144;
squeal_samples[1448]=10311;
squeal_samples[1449]=13472;
squeal_samples[1450]=16494;
squeal_samples[1451]=19392;
squeal_samples[1452]=22160;
squeal_samples[1453]=24814;
squeal_samples[1454]=27352;
squeal_samples[1455]=29773;
squeal_samples[1456]=32092;
squeal_samples[1457]=34306;
squeal_samples[1458]=36428;
squeal_samples[1459]=38448;
squeal_samples[1460]=40383;
squeal_samples[1461]=42229;
squeal_samples[1462]=43996;
squeal_samples[1463]=45685;
squeal_samples[1464]=47292;
squeal_samples[1465]=48836;
squeal_samples[1466]=50306;
squeal_samples[1467]=49883;
squeal_samples[1468]=45090;
squeal_samples[1469]=40426;
squeal_samples[1470]=36051;
squeal_samples[1471]=31961;
squeal_samples[1472]=28138;
squeal_samples[1473]=24554;
squeal_samples[1474]=21202;
squeal_samples[1475]=18071;
squeal_samples[1476]=15140;
squeal_samples[1477]=12399;
squeal_samples[1478]=9837;
squeal_samples[1479]=8139;
squeal_samples[1480]=10703;
squeal_samples[1481]=13841;
squeal_samples[1482]=16848;
squeal_samples[1483]=19729;
squeal_samples[1484]=22489;
squeal_samples[1485]=25127;
squeal_samples[1486]=27647;
squeal_samples[1487]=30060;
squeal_samples[1488]=32359;
squeal_samples[1489]=34559;
squeal_samples[1490]=36675;
squeal_samples[1491]=38679;
squeal_samples[1492]=40609;
squeal_samples[1493]=42442;
squeal_samples[1494]=44197;
squeal_samples[1495]=45875;
squeal_samples[1496]=47477;
squeal_samples[1497]=49011;
squeal_samples[1498]=50474;
squeal_samples[1499]=49380;
squeal_samples[1500]=44480;
squeal_samples[1501]=39847;
squeal_samples[1502]=35509;
squeal_samples[1503]=31457;
squeal_samples[1504]=27661;
squeal_samples[1505]=24113;
squeal_samples[1506]=20789;
squeal_samples[1507]=17678;
squeal_samples[1508]=14780;
squeal_samples[1509]=12055;
squeal_samples[1510]=9517;
squeal_samples[1511]=8234;
squeal_samples[1512]=11092;
squeal_samples[1513]=14208;
squeal_samples[1514]=17206;
squeal_samples[1515]=20067;
squeal_samples[1516]=22815;
squeal_samples[1517]=25432;
squeal_samples[1518]=27945;
squeal_samples[1519]=30335;
squeal_samples[1520]=32627;
squeal_samples[1521]=34821;
squeal_samples[1522]=36912;
squeal_samples[1523]=38917;
squeal_samples[1524]=40823;
squeal_samples[1525]=42658;
squeal_samples[1526]=44397;
squeal_samples[1527]=46072;
squeal_samples[1528]=47657;
squeal_samples[1529]=49186;
squeal_samples[1530]=50639;
squeal_samples[1531]=48787;
squeal_samples[1532]=43869;
squeal_samples[1533]=39279;
squeal_samples[1534]=34978;
squeal_samples[1535]=30952;
squeal_samples[1536]=27196;
squeal_samples[1537]=23669;
squeal_samples[1538]=20374;
squeal_samples[1539]=17293;
squeal_samples[1540]=14412;
squeal_samples[1541]=11713;
squeal_samples[1542]=9199;
squeal_samples[1543]=8412;
squeal_samples[1544]=11475;
squeal_samples[1545]=14579;
squeal_samples[1546]=17553;
squeal_samples[1547]=20406;
squeal_samples[1548]=23131;
squeal_samples[1549]=25741;
squeal_samples[1550]=28237;
squeal_samples[1551]=30613;
squeal_samples[1552]=32901;
squeal_samples[1553]=35069;
squeal_samples[1554]=37162;
squeal_samples[1555]=39141;
squeal_samples[1556]=41052;
squeal_samples[1557]=42861;
squeal_samples[1558]=44602;
squeal_samples[1559]=46257;
squeal_samples[1560]=47844;
squeal_samples[1561]=49354;
squeal_samples[1562]=50757;
squeal_samples[1563]=48134;
squeal_samples[1564]=43269;
squeal_samples[1565]=38710;
squeal_samples[1566]=34450;
squeal_samples[1567]=30457;
squeal_samples[1568]=26726;
squeal_samples[1569]=23236;
squeal_samples[1570]=19962;
squeal_samples[1571]=16916;
squeal_samples[1572]=14052;
squeal_samples[1573]=11384;
squeal_samples[1574]=8880;
squeal_samples[1575]=8679;
squeal_samples[1576]=11859;
squeal_samples[1577]=14947;
squeal_samples[1578]=17904;
squeal_samples[1579]=20742;
squeal_samples[1580]=23451;
squeal_samples[1581]=26044;
squeal_samples[1582]=28527;
squeal_samples[1583]=30892;
squeal_samples[1584]=33161;
squeal_samples[1585]=35329;
squeal_samples[1586]=37400;
squeal_samples[1587]=39376;
squeal_samples[1588]=41267;
squeal_samples[1589]=43072;
squeal_samples[1590]=44802;
squeal_samples[1591]=46445;
squeal_samples[1592]=48023;
squeal_samples[1593]=49528;
squeal_samples[1594]=50766;
squeal_samples[1595]=47498;
squeal_samples[1596]=42674;
squeal_samples[1597]=38150;
squeal_samples[1598]=33924;
squeal_samples[1599]=29965;
squeal_samples[1600]=26271;
squeal_samples[1601]=22804;
squeal_samples[1602]=19561;
squeal_samples[1603]=16532;
squeal_samples[1604]=13695;
squeal_samples[1605]=11051;
squeal_samples[1606]=8570;
squeal_samples[1607]=9029;
squeal_samples[1608]=12242;
squeal_samples[1609]=15311;
squeal_samples[1610]=18261;
squeal_samples[1611]=21077;
squeal_samples[1612]=23768;
squeal_samples[1613]=26198;
squeal_samples[1614]=28513;
squeal_samples[1615]=30881;
squeal_samples[1616]=33150;
squeal_samples[1617]=35315;
squeal_samples[1618]=37390;
squeal_samples[1619]=39363;
squeal_samples[1620]=41256;
squeal_samples[1621]=43060;
squeal_samples[1622]=44790;
squeal_samples[1623]=46433;
squeal_samples[1624]=48013;
squeal_samples[1625]=49513;
squeal_samples[1626]=50758;
squeal_samples[1627]=47484;
squeal_samples[1628]=42662;
squeal_samples[1629]=38141;
squeal_samples[1630]=33910;
squeal_samples[1631]=29953;
squeal_samples[1632]=26261;
squeal_samples[1633]=22789;
squeal_samples[1634]=19554;
squeal_samples[1635]=16517;
squeal_samples[1636]=13687;
squeal_samples[1637]=11034;
squeal_samples[1638]=8563;
squeal_samples[1639]=9015;
squeal_samples[1640]=12231;
squeal_samples[1641]=15301;
squeal_samples[1642]=18248;
squeal_samples[1643]=21064;
squeal_samples[1644]=23760;
squeal_samples[1645]=26339;
squeal_samples[1646]=28811;
squeal_samples[1647]=31153;
squeal_samples[1648]=33418;
squeal_samples[1649]=35569;
squeal_samples[1650]=37628;
squeal_samples[1651]=39591;
squeal_samples[1652]=41478;
squeal_samples[1653]=43265;
squeal_samples[1654]=44987;
squeal_samples[1655]=46622;
squeal_samples[1656]=48196;
squeal_samples[1657]=49689;
squeal_samples[1658]=50664;
squeal_samples[1659]=46852;
squeal_samples[1660]=42073;
squeal_samples[1661]=37582;
squeal_samples[1662]=33390;
squeal_samples[1663]=29472;
squeal_samples[1664]=25799;
squeal_samples[1665]=22365;
squeal_samples[1666]=19147;
squeal_samples[1667]=16145;
squeal_samples[1668]=13332;
squeal_samples[1669]=10704;
squeal_samples[1670]=8292;
squeal_samples[1671]=9415;
squeal_samples[1672]=12610;
squeal_samples[1673]=15664;
squeal_samples[1674]=18596;
squeal_samples[1675]=21394;
squeal_samples[1676]=24080;
squeal_samples[1677]=26638;
squeal_samples[1678]=29096;
squeal_samples[1679]=31433;
squeal_samples[1680]=33675;
squeal_samples[1681]=35821;
squeal_samples[1682]=37863;
squeal_samples[1683]=39828;
squeal_samples[1684]=41691;
squeal_samples[1685]=43480;
squeal_samples[1686]=45184;
squeal_samples[1687]=46813;
squeal_samples[1688]=48374;
squeal_samples[1689]=49858;
squeal_samples[1690]=50824;
squeal_samples[1691]=47009;
squeal_samples[1692]=42206;
squeal_samples[1693]=37720;
squeal_samples[1694]=33508;
squeal_samples[1695]=29589;
squeal_samples[1696]=25902;
squeal_samples[1697]=22461;
squeal_samples[1698]=19240;
squeal_samples[1699]=16226;
squeal_samples[1700]=13412;
squeal_samples[1701]=10775;
squeal_samples[1702]=8363;
squeal_samples[1703]=9479;
squeal_samples[1704]=12669;
squeal_samples[1705]=15719;
squeal_samples[1706]=18649;
squeal_samples[1707]=21444;
squeal_samples[1708]=24127;
squeal_samples[1709]=26689;
squeal_samples[1710]=29136;
squeal_samples[1711]=31479;
squeal_samples[1712]=33717;
squeal_samples[1713]=35859;
squeal_samples[1714]=37902;
squeal_samples[1715]=39858;
squeal_samples[1716]=41726;
squeal_samples[1717]=43506;
squeal_samples[1718]=45211;
squeal_samples[1719]=46841;
squeal_samples[1720]=48396;
squeal_samples[1721]=49886;
squeal_samples[1722]=50487;
squeal_samples[1723]=46247;
squeal_samples[1724]=41496;
squeal_samples[1725]=37051;
squeal_samples[1726]=32885;
squeal_samples[1727]=29001;
squeal_samples[1728]=25354;
squeal_samples[1729]=21945;
squeal_samples[1730]=18757;
squeal_samples[1731]=15775;
squeal_samples[1732]=12988;
squeal_samples[1733]=10386;
squeal_samples[1734]=8120;
squeal_samples[1735]=9816;
squeal_samples[1736]=12985;
squeal_samples[1737]=16032;
squeal_samples[1738]=18939;
squeal_samples[1739]=21730;
squeal_samples[1740]=24390;
squeal_samples[1741]=26948;
squeal_samples[1742]=29378;
squeal_samples[1743]=31712;
squeal_samples[1744]=33935;
squeal_samples[1745]=36069;
squeal_samples[1746]=38105;
squeal_samples[1747]=40048;
squeal_samples[1748]=41904;
squeal_samples[1749]=43679;
squeal_samples[1750]=45375;
squeal_samples[1751]=46997;
squeal_samples[1752]=48550;
squeal_samples[1753]=50025;
squeal_samples[1754]=50625;
squeal_samples[1755]=46368;
squeal_samples[1756]=41615;
squeal_samples[1757]=37154;
squeal_samples[1758]=32994;
squeal_samples[1759]=29088;
squeal_samples[1760]=25444;
squeal_samples[1761]=22025;
squeal_samples[1762]=18834;
squeal_samples[1763]=15845;
squeal_samples[1764]=13053;
squeal_samples[1765]=10445;
squeal_samples[1766]=8177;
squeal_samples[1767]=9867;
squeal_samples[1768]=13036;
squeal_samples[1769]=16074;
squeal_samples[1770]=18985;
squeal_samples[1771]=21771;
squeal_samples[1772]=24431;
squeal_samples[1773]=26981;
squeal_samples[1774]=29420;
squeal_samples[1775]=31744;
squeal_samples[1776]=33967;
squeal_samples[1777]=36098;
squeal_samples[1778]=38130;
squeal_samples[1779]=40076;
squeal_samples[1780]=41930;
squeal_samples[1781]=43704;
squeal_samples[1782]=45394;
squeal_samples[1783]=47016;
squeal_samples[1784]=48564;
squeal_samples[1785]=50042;
squeal_samples[1786]=50641;
squeal_samples[1787]=46387;
squeal_samples[1788]=41627;
squeal_samples[1789]=37171;
squeal_samples[1790]=32991;
squeal_samples[1791]=29109;
squeal_samples[1792]=25446;
squeal_samples[1793]=22043;
squeal_samples[1794]=18835;
squeal_samples[1795]=15853;
squeal_samples[1796]=13057;
squeal_samples[1797]=10448;
squeal_samples[1798]=8173;
squeal_samples[1799]=9871;
squeal_samples[1800]=13034;
squeal_samples[1801]=16075;
squeal_samples[1802]=18986;
squeal_samples[1803]=21768;
squeal_samples[1804]=24433;
squeal_samples[1805]=26982;
squeal_samples[1806]=29414;
squeal_samples[1807]=31739;
squeal_samples[1808]=33967;
squeal_samples[1809]=36097;
squeal_samples[1810]=38127;
squeal_samples[1811]=40069;
squeal_samples[1812]=41926;
squeal_samples[1813]=43699;
squeal_samples[1814]=45387;
squeal_samples[1815]=47014;
squeal_samples[1816]=48555;
squeal_samples[1817]=50039;
squeal_samples[1818]=50636;
squeal_samples[1819]=46381;
squeal_samples[1820]=41618;
squeal_samples[1821]=37163;
squeal_samples[1822]=32989;
squeal_samples[1823]=29100;
squeal_samples[1824]=25441;
squeal_samples[1825]=22026;
squeal_samples[1826]=18835;
squeal_samples[1827]=15844;
squeal_samples[1828]=13051;
squeal_samples[1829]=10432;
squeal_samples[1830]=8173;
squeal_samples[1831]=9860;
squeal_samples[1832]=13029;
squeal_samples[1833]=16061;
squeal_samples[1834]=18976;
squeal_samples[1835]=21759;
squeal_samples[1836]=24426;
squeal_samples[1837]=26972;
squeal_samples[1838]=29409;
squeal_samples[1839]=31733;
squeal_samples[1840]=33958;
squeal_samples[1841]=36086;
squeal_samples[1842]=38116;
squeal_samples[1843]=40058;
squeal_samples[1844]=41917;
squeal_samples[1845]=43691;
squeal_samples[1846]=45386;
squeal_samples[1847]=47004;
squeal_samples[1848]=48548;
squeal_samples[1849]=50028;
squeal_samples[1850]=50623;
squeal_samples[1851]=46374;
squeal_samples[1852]=41609;
squeal_samples[1853]=37155;
squeal_samples[1854]=32978;
squeal_samples[1855]=29089;
squeal_samples[1856]=25430;
squeal_samples[1857]=22018;
squeal_samples[1858]=18821;
squeal_samples[1859]=15837;
squeal_samples[1860]=13037;
squeal_samples[1861]=10428;
squeal_samples[1862]=8163;
squeal_samples[1863]=9851;
squeal_samples[1864]=13021;
squeal_samples[1865]=16058;
squeal_samples[1866]=18963;
squeal_samples[1867]=21751;
squeal_samples[1868]=24414;
squeal_samples[1869]=26963;
squeal_samples[1870]=29397;
squeal_samples[1871]=31722;
squeal_samples[1872]=33949;
squeal_samples[1873]=36073;
squeal_samples[1874]=38108;
squeal_samples[1875]=40046;
squeal_samples[1876]=41907;
squeal_samples[1877]=43679;
squeal_samples[1878]=45377;
squeal_samples[1879]=46993;
squeal_samples[1880]=48538;
squeal_samples[1881]=50017;
squeal_samples[1882]=50612;
squeal_samples[1883]=46363;
squeal_samples[1884]=41601;
squeal_samples[1885]=37141;
squeal_samples[1886]=32972;
squeal_samples[1887]=29073;
squeal_samples[1888]=25424;
squeal_samples[1889]=22003;
squeal_samples[1890]=18814;
squeal_samples[1891]=15823;
squeal_samples[1892]=13030;
squeal_samples[1893]=10415;
squeal_samples[1894]=8153;
squeal_samples[1895]=9840;
squeal_samples[1896]=13010;
squeal_samples[1897]=16049;
squeal_samples[1898]=18952;
squeal_samples[1899]=21738;
squeal_samples[1900]=24408;
squeal_samples[1901]=26947;
squeal_samples[1902]=29392;
squeal_samples[1903]=31708;
squeal_samples[1904]=33939;
squeal_samples[1905]=36064;
squeal_samples[1906]=38095;
squeal_samples[1907]=40038;
squeal_samples[1908]=41894;
squeal_samples[1909]=43671;
squeal_samples[1910]=45364;
squeal_samples[1911]=46984;
squeal_samples[1912]=48525;
squeal_samples[1913]=50009;
squeal_samples[1914]=50600;
squeal_samples[1915]=46353;
squeal_samples[1916]=41589;
squeal_samples[1917]=37132;
squeal_samples[1918]=32960;
squeal_samples[1919]=29063;
squeal_samples[1920]=25414;
squeal_samples[1921]=21991;
squeal_samples[1922]=18805;
squeal_samples[1923]=15813;
squeal_samples[1924]=13017;
squeal_samples[1925]=10407;
squeal_samples[1926]=8140;
squeal_samples[1927]=9831;
squeal_samples[1928]=12999;
squeal_samples[1929]=16039;
squeal_samples[1930]=18941;
squeal_samples[1931]=21728;
squeal_samples[1932]=24396;
squeal_samples[1933]=26937;
squeal_samples[1934]=29381;
squeal_samples[1935]=31699;
squeal_samples[1936]=33927;
squeal_samples[1937]=36053;
squeal_samples[1938]=38085;
squeal_samples[1939]=40026;
squeal_samples[1940]=41887;
squeal_samples[1941]=43657;
squeal_samples[1942]=45354;
squeal_samples[1943]=46974;
squeal_samples[1944]=48515;
squeal_samples[1945]=49996;
squeal_samples[1946]=50594;
squeal_samples[1947]=46337;
squeal_samples[1948]=41583;
squeal_samples[1949]=37119;
squeal_samples[1950]=32949;
squeal_samples[1951]=29055;
squeal_samples[1952]=25400;
squeal_samples[1953]=21983;
squeal_samples[1954]=18793;
squeal_samples[1955]=15802;
squeal_samples[1956]=13007;
squeal_samples[1957]=10396;
squeal_samples[1958]=8130;
squeal_samples[1959]=9819;
squeal_samples[1960]=12990;
squeal_samples[1961]=16025;
squeal_samples[1962]=18934;
squeal_samples[1963]=21716;
squeal_samples[1964]=24384;
squeal_samples[1965]=26929;
squeal_samples[1966]=29366;
squeal_samples[1967]=31693;
squeal_samples[1968]=33912;
squeal_samples[1969]=36046;
squeal_samples[1970]=38071;
squeal_samples[1971]=40018;
squeal_samples[1972]=41874;
squeal_samples[1973]=43646;
squeal_samples[1974]=45346;
squeal_samples[1975]=46960;
squeal_samples[1976]=48506;
squeal_samples[1977]=49986;
squeal_samples[1978]=50580;
squeal_samples[1979]=46330;
squeal_samples[1980]=41570;
squeal_samples[1981]=37108;
squeal_samples[1982]=32939;
squeal_samples[1983]=29044;
squeal_samples[1984]=25389;
squeal_samples[1985]=21974;
squeal_samples[1986]=18780;
squeal_samples[1987]=15791;
squeal_samples[1988]=12998;
squeal_samples[1989]=10383;
squeal_samples[1990]=8121;
squeal_samples[1991]=9808;
squeal_samples[1992]=12978;
squeal_samples[1993]=16016;
squeal_samples[1994]=18921;
squeal_samples[1995]=21706;
squeal_samples[1996]=24373;
squeal_samples[1997]=26918;
squeal_samples[1998]=29357;
squeal_samples[1999]=31679;
squeal_samples[2000]=33904;
squeal_samples[2001]=36034;
squeal_samples[2002]=38060;
squeal_samples[2003]=40008;
squeal_samples[2004]=41862;
squeal_samples[2005]=43636;
squeal_samples[2006]=45336;
squeal_samples[2007]=46948;
squeal_samples[2008]=48496;
squeal_samples[2009]=49973;
squeal_samples[2010]=50572;
squeal_samples[2011]=46316;
squeal_samples[2012]=41562;
squeal_samples[2013]=37096;
squeal_samples[2014]=32928;
squeal_samples[2015]=29032;
squeal_samples[2016]=25380;
squeal_samples[2017]=21960;
squeal_samples[2018]=18773;
squeal_samples[2019]=15778;
squeal_samples[2020]=12986;
squeal_samples[2021]=10375;
squeal_samples[2022]=8108;
squeal_samples[2023]=9796;
squeal_samples[2024]=12971;
squeal_samples[2025]=16000;
squeal_samples[2026]=18914;
squeal_samples[2027]=21693;
squeal_samples[2028]=24362;
squeal_samples[2029]=26908;
squeal_samples[2030]=29345;
squeal_samples[2031]=31667;
squeal_samples[2032]=33896;
squeal_samples[2033]=36019;
squeal_samples[2034]=38053;
squeal_samples[2035]=39993;
squeal_samples[2036]=41852;
squeal_samples[2037]=43627;
squeal_samples[2038]=45322;
squeal_samples[2039]=46938;
squeal_samples[2040]=48484;
squeal_samples[2041]=49962;
squeal_samples[2042]=50917;
squeal_samples[2043]=47086;
squeal_samples[2044]=42274;
squeal_samples[2045]=37772;
squeal_samples[2046]=33557;
squeal_samples[2047]=29618;
squeal_samples[2048]=25928;
squeal_samples[2049]=22477;
squeal_samples[2050]=19246;
squeal_samples[2051]=16230;
squeal_samples[2052]=13397;
squeal_samples[2053]=10766;
squeal_samples[2054]=8331;
squeal_samples[2055]=9459;
squeal_samples[2056]=12633;
squeal_samples[2057]=15685;
squeal_samples[2058]=18604;
squeal_samples[2059]=21408;
squeal_samples[2060]=24081;
squeal_samples[2061]=26639;
squeal_samples[2062]=29091;
squeal_samples[2063]=31422;
squeal_samples[2064]=33660;
squeal_samples[2065]=35801;
squeal_samples[2066]=37837;
squeal_samples[2067]=39790;
squeal_samples[2068]=41653;
squeal_samples[2069]=43439;
squeal_samples[2070]=45134;
squeal_samples[2071]=46769;
squeal_samples[2072]=48316;
squeal_samples[2073]=49809;
squeal_samples[2074]=50762;
squeal_samples[2075]=46945;
squeal_samples[2076]=42138;
squeal_samples[2077]=37647;
squeal_samples[2078]=33437;
squeal_samples[2079]=29506;
squeal_samples[2080]=25822;
squeal_samples[2081]=22375;
squeal_samples[2082]=19153;
squeal_samples[2083]=16141;
squeal_samples[2084]=13321;
squeal_samples[2085]=10682;
squeal_samples[2086]=8269;
squeal_samples[2087]=9379;
squeal_samples[2088]=12569;
squeal_samples[2089]=15615;
squeal_samples[2090]=18547;
squeal_samples[2091]=21342;
squeal_samples[2092]=24019;
squeal_samples[2093]=26580;
squeal_samples[2094]=29036;
squeal_samples[2095]=31368;
squeal_samples[2096]=33606;
squeal_samples[2097]=35744;
squeal_samples[2098]=37789;
squeal_samples[2099]=39746;
squeal_samples[2100]=41610;
squeal_samples[2101]=43393;
squeal_samples[2102]=45098;
squeal_samples[2103]=46721;
squeal_samples[2104]=48282;
squeal_samples[2105]=49766;
squeal_samples[2106]=50981;
squeal_samples[2107]=47693;
squeal_samples[2108]=42838;
squeal_samples[2109]=38301;
squeal_samples[2110]=34046;
squeal_samples[2111]=30078;
squeal_samples[2112]=26358;
squeal_samples[2113]=22874;
squeal_samples[2114]=19622;
squeal_samples[2115]=16572;
squeal_samples[2116]=13728;
squeal_samples[2117]=11063;
squeal_samples[2118]=8576;
squeal_samples[2119]=9022;
squeal_samples[2120]=12231;
squeal_samples[2121]=15286;
squeal_samples[2122]=18236;
squeal_samples[2123]=21037;
squeal_samples[2124]=23735;
squeal_samples[2125]=26301;
squeal_samples[2126]=28769;
squeal_samples[2127]=31114;
squeal_samples[2128]=33365;
squeal_samples[2129]=35516;
squeal_samples[2130]=37566;
squeal_samples[2131]=39533;
squeal_samples[2132]=41403;
squeal_samples[2133]=43198;
squeal_samples[2134]=44905;
squeal_samples[2135]=46544;
squeal_samples[2136]=48104;
squeal_samples[2137]=49604;
squeal_samples[2138]=50979;
squeal_samples[2139]=48338;
squeal_samples[2140]=43445;
squeal_samples[2141]=38858;
squeal_samples[2142]=34580;
squeal_samples[2143]=30560;
squeal_samples[2144]=26817;
squeal_samples[2145]=23301;
squeal_samples[2146]=20022;
squeal_samples[2147]=16947;
squeal_samples[2148]=14075;
squeal_samples[2149]=11384;
squeal_samples[2150]=8878;
squeal_samples[2151]=8659;
squeal_samples[2152]=11830;
squeal_samples[2153]=14916;
squeal_samples[2154]=17864;
squeal_samples[2155]=20696;
squeal_samples[2156]=23398;
squeal_samples[2157]=25988;
squeal_samples[2158]=28465;
squeal_samples[2159]=30822;
squeal_samples[2160]=33085;
squeal_samples[2161]=35247;
squeal_samples[2162]=37312;
squeal_samples[2163]=39287;
squeal_samples[2164]=41170;
squeal_samples[2165]=42973;
squeal_samples[2166]=44694;
squeal_samples[2167]=46340;
squeal_samples[2168]=47910;
squeal_samples[2169]=49412;
squeal_samples[2170]=50847;
squeal_samples[2171]=48964;
squeal_samples[2172]=44028;
squeal_samples[2173]=39409;
squeal_samples[2174]=35087;
squeal_samples[2175]=31046;
squeal_samples[2176]=27262;
squeal_samples[2177]=23729;
squeal_samples[2178]=20407;
squeal_samples[2179]=17316;
squeal_samples[2180]=14412;
squeal_samples[2181]=11706;
squeal_samples[2182]=9170;
squeal_samples[2183]=8376;
squeal_samples[2184]=11427;
squeal_samples[2185]=14523;
squeal_samples[2186]=17496;
squeal_samples[2187]=20340;
squeal_samples[2188]=23062;
squeal_samples[2189]=25660;
squeal_samples[2190]=28149;
squeal_samples[2191]=30524;
squeal_samples[2192]=32800;
squeal_samples[2193]=34971;
squeal_samples[2194]=37049;
squeal_samples[2195]=39032;
squeal_samples[2196]=40928;
squeal_samples[2197]=42741;
squeal_samples[2198]=44470;
squeal_samples[2199]=46126;
squeal_samples[2200]=47711;
squeal_samples[2201]=49210;
squeal_samples[2202]=50665;
squeal_samples[2203]=49544;
squeal_samples[2204]=44618;
squeal_samples[2205]=39965;
squeal_samples[2206]=35600;
squeal_samples[2207]=31522;
squeal_samples[2208]=27710;
squeal_samples[2209]=24141;
squeal_samples[2210]=20803;
squeal_samples[2211]=17674;
squeal_samples[2212]=14751;
squeal_samples[2213]=12017;
squeal_samples[2214]=9471;
squeal_samples[2215]=8172;
squeal_samples[2216]=11019;
squeal_samples[2217]=14137;
squeal_samples[2218]=17118;
squeal_samples[2219]=19977;
squeal_samples[2220]=22712;
squeal_samples[2221]=25329;
squeal_samples[2222]=27832;
squeal_samples[2223]=30221;
squeal_samples[2224]=32504;
squeal_samples[2225]=34695;
squeal_samples[2226]=36780;
squeal_samples[2227]=38782;
squeal_samples[2228]=40684;
squeal_samples[2229]=42505;
squeal_samples[2230]=44246;
squeal_samples[2231]=45910;
squeal_samples[2232]=47500;
squeal_samples[2233]=49017;
squeal_samples[2234]=50471;
squeal_samples[2235]=50021;
squeal_samples[2236]=45211;
squeal_samples[2237]=40515;
squeal_samples[2238]=36123;
squeal_samples[2239]=32003;
squeal_samples[2240]=28166;
squeal_samples[2241]=24564;
squeal_samples[2242]=21191;
squeal_samples[2243]=18042;
squeal_samples[2244]=15099;
squeal_samples[2245]=12342;
squeal_samples[2246]=9768;
squeal_samples[2247]=8059;
squeal_samples[2248]=10606;
squeal_samples[2249]=13743;
squeal_samples[2250]=16740;
squeal_samples[2251]=19619;
squeal_samples[2252]=22363;
squeal_samples[2253]=24996;
squeal_samples[2254]=27517;
squeal_samples[2255]=29915;
squeal_samples[2256]=32216;
squeal_samples[2257]=34416;
squeal_samples[2258]=36514;
squeal_samples[2259]=38519;
squeal_samples[2260]=40440;
squeal_samples[2261]=42269;
squeal_samples[2262]=44023;
squeal_samples[2263]=45696;
squeal_samples[2264]=47292;
squeal_samples[2265]=48822;
squeal_samples[2266]=50276;
squeal_samples[2267]=50398;
squeal_samples[2268]=45805;
squeal_samples[2269]=41076;
squeal_samples[2270]=36641;
squeal_samples[2271]=32491;
squeal_samples[2272]=28622;
squeal_samples[2273]=24983;
squeal_samples[2274]=21596;
squeal_samples[2275]=18413;
squeal_samples[2276]=15440;
squeal_samples[2277]=12663;
squeal_samples[2278]=10063;
squeal_samples[2279]=8032;
squeal_samples[2280]=10193;
squeal_samples[2281]=13347;
squeal_samples[2282]=16364;
squeal_samples[2283]=19248;
squeal_samples[2284]=22018;
squeal_samples[2285]=24662;
squeal_samples[2286]=27196;
squeal_samples[2287]=29614;
squeal_samples[2288]=31924;
squeal_samples[2289]=34130;
squeal_samples[2290]=36243;
squeal_samples[2291]=38261;
squeal_samples[2292]=40196;
squeal_samples[2293]=42032;
squeal_samples[2294]=43797;
squeal_samples[2295]=45473;
squeal_samples[2296]=47088;
squeal_samples[2297]=48622;
squeal_samples[2298]=50092;
squeal_samples[2299]=50672;
squeal_samples[2300]=46408;
squeal_samples[2301]=41633;
squeal_samples[2302]=37167;
squeal_samples[2303]=32984;
squeal_samples[2304]=29076;
squeal_samples[2305]=25413;
squeal_samples[2306]=21993;
squeal_samples[2307]=18790;
squeal_samples[2308]=15787;
squeal_samples[2309]=12992;
squeal_samples[2310]=10364;
squeal_samples[2311]=8096;
squeal_samples[2312]=9779;
squeal_samples[2313]=12943;
squeal_samples[2314]=15980;
squeal_samples[2315]=18888;
squeal_samples[2316]=21663;
squeal_samples[2317]=24329;
squeal_samples[2318]=26871;
squeal_samples[2319]=29304;
squeal_samples[2320]=31625;
squeal_samples[2321]=33844;
squeal_samples[2322]=35977;
squeal_samples[2323]=38005;
squeal_samples[2324]=39941;
squeal_samples[2325]=41798;
squeal_samples[2326]=43566;
squeal_samples[2327]=45260;
squeal_samples[2328]=46877;
squeal_samples[2329]=48419;
squeal_samples[2330]=49902;
squeal_samples[2331]=50847;
squeal_samples[2332]=47018;
squeal_samples[2333]=42200;
squeal_samples[2334]=37699;
squeal_samples[2335]=33477;
squeal_samples[2336]=29539;
squeal_samples[2337]=25849;
squeal_samples[2338]=22390;
squeal_samples[2339]=19166;
squeal_samples[2340]=16138;
squeal_samples[2341]=13320;
squeal_samples[2342]=10674;
squeal_samples[2343]=8252;
squeal_samples[2344]=9363;
squeal_samples[2345]=12547;
squeal_samples[2346]=15591;
squeal_samples[2347]=18516;
squeal_samples[2348]=21312;
squeal_samples[2349]=23987;
squeal_samples[2350]=26546;
squeal_samples[2351]=28993;
squeal_samples[2352]=31327;
squeal_samples[2353]=33565;
squeal_samples[2354]=35699;
squeal_samples[2355]=37747;
squeal_samples[2356]=39688;
squeal_samples[2357]=41562;
squeal_samples[2358]=43338;
squeal_samples[2359]=45040;
squeal_samples[2360]=46662;
squeal_samples[2361]=48220;
squeal_samples[2362]=49701;
squeal_samples[2363]=50917;
squeal_samples[2364]=47632;
squeal_samples[2365]=42771;
squeal_samples[2366]=38232;
squeal_samples[2367]=33980;
squeal_samples[2368]=29999;
squeal_samples[2369]=26287;
squeal_samples[2370]=22797;
squeal_samples[2371]=19541;
squeal_samples[2372]=16493;
squeal_samples[2373]=13647;
squeal_samples[2374]=10984;
squeal_samples[2375]=8493;
squeal_samples[2376]=8945;
squeal_samples[2377]=12140;
squeal_samples[2378]=15206;
squeal_samples[2379]=18144;
squeal_samples[2380]=20956;
squeal_samples[2381]=23646;
squeal_samples[2382]=26216;
squeal_samples[2383]=28683;
squeal_samples[2384]=31026;
squeal_samples[2385]=33274;
squeal_samples[2386]=35425;
squeal_samples[2387]=37479;
squeal_samples[2388]=39441;
squeal_samples[2389]=41318;
squeal_samples[2390]=43103;
squeal_samples[2391]=44824;
squeal_samples[2392]=46451;
squeal_samples[2393]=48018;
squeal_samples[2394]=49507;
squeal_samples[2395]=50891;
squeal_samples[2396]=48246;
squeal_samples[2397]=43349;
squeal_samples[2398]=38771;
squeal_samples[2399]=34482;
squeal_samples[2400]=30473;
squeal_samples[2401]=26722;
squeal_samples[2402]=23210;
squeal_samples[2403]=19923;
squeal_samples[2404]=16851;
squeal_samples[2405]=13975;
squeal_samples[2406]=11293;
squeal_samples[2407]=8780;
squeal_samples[2408]=8566;
squeal_samples[2409]=11739;
squeal_samples[2410]=14815;
squeal_samples[2411]=17775;
squeal_samples[2412]=20595;
squeal_samples[2413]=23307;
squeal_samples[2414]=25889;
squeal_samples[2415]=28366;
squeal_samples[2416]=30725;
squeal_samples[2417]=32992;
squeal_samples[2418]=35148;
squeal_samples[2419]=37213;
squeal_samples[2420]=39189;
squeal_samples[2421]=41071;
squeal_samples[2422]=42875;
squeal_samples[2423]=44595;
squeal_samples[2424]=46241;
squeal_samples[2425]=47811;
squeal_samples[2426]=49312;
squeal_samples[2427]=50749;
squeal_samples[2428]=49620;
squeal_samples[2429]=44685;
squeal_samples[2430]=40016;
squeal_samples[2431]=35650;
squeal_samples[2432]=31565;
squeal_samples[2433]=27742;
squeal_samples[2434]=24164;
squeal_samples[2435]=20816;
squeal_samples[2436]=17687;
squeal_samples[2437]=14752;
squeal_samples[2438]=12022;
squeal_samples[2439]=9454;
squeal_samples[2440]=8160;
squeal_samples[2441]=11004;
squeal_samples[2442]=14117;
squeal_samples[2443]=17094;
squeal_samples[2444]=19956;
squeal_samples[2445]=22683;
squeal_samples[2446]=25302;
squeal_samples[2447]=27800;
squeal_samples[2448]=30184;
squeal_samples[2449]=32475;
squeal_samples[2450]=34652;
squeal_samples[2451]=36738;
squeal_samples[2452]=38738;
squeal_samples[2453]=40637;
squeal_samples[2454]=42463;
squeal_samples[2455]=44195;
squeal_samples[2456]=45859;
squeal_samples[2457]=47445;
squeal_samples[2458]=48967;
squeal_samples[2459]=50413;
squeal_samples[2460]=50522;
squeal_samples[2461]=45915;
squeal_samples[2462]=41172;
squeal_samples[2463]=36728;
squeal_samples[2464]=32573;
squeal_samples[2465]=28686;
squeal_samples[2466]=25045;
squeal_samples[2467]=21642;
squeal_samples[2468]=18452;
squeal_samples[2469]=15477;
squeal_samples[2470]=12691;
squeal_samples[2471]=10084;
squeal_samples[2472]=8047;
squeal_samples[2473]=10204;
squeal_samples[2474]=13353;
squeal_samples[2475]=16362;
squeal_samples[2476]=19249;
squeal_samples[2477]=22016;
squeal_samples[2478]=24652;
squeal_samples[2479]=27183;
squeal_samples[2480]=29600;
squeal_samples[2481]=31903;
squeal_samples[2482]=34117;
squeal_samples[2483]=36218;
squeal_samples[2484]=38241;
squeal_samples[2485]=40165;
squeal_samples[2486]=42009;
squeal_samples[2487]=43763;
squeal_samples[2488]=45446;
squeal_samples[2489]=47050;
squeal_samples[2490]=48585;
squeal_samples[2491]=50052;
squeal_samples[2492]=50991;
squeal_samples[2493]=47147;
squeal_samples[2494]=42323;
squeal_samples[2495]=37800;
squeal_samples[2496]=33577;
squeal_samples[2497]=29626;
squeal_samples[2498]=25925;
squeal_samples[2499]=22459;
squeal_samples[2500]=19221;
squeal_samples[2501]=16193;
squeal_samples[2502]=13354;
squeal_samples[2503]=10710;
squeal_samples[2504]=8278;
squeal_samples[2505]=9387;
squeal_samples[2506]=12567;
squeal_samples[2507]=15609;
squeal_samples[2508]=18533;
squeal_samples[2509]=21321;
squeal_samples[2510]=23996;
squeal_samples[2511]=26550;
squeal_samples[2512]=28993;
squeal_samples[2513]=31324;
squeal_samples[2514]=33557;
squeal_samples[2515]=35692;
squeal_samples[2516]=37733;
squeal_samples[2517]=39680;
squeal_samples[2518]=41544;
squeal_samples[2519]=43318;
squeal_samples[2520]=45017;
squeal_samples[2521]=46643;
squeal_samples[2522]=48194;
squeal_samples[2523]=49682;
squeal_samples[2524]=51047;
squeal_samples[2525]=48396;
squeal_samples[2526]=43487;
squeal_samples[2527]=38891;
squeal_samples[2528]=34595;
squeal_samples[2529]=30569;
squeal_samples[2530]=26815;
squeal_samples[2531]=23289;
squeal_samples[2532]=20001;
squeal_samples[2533]=16912;
squeal_samples[2534]=14042;
squeal_samples[2535]=11340;
squeal_samples[2536]=8827;
squeal_samples[2537]=8601;
squeal_samples[2538]=11771;
squeal_samples[2539]=14847;
squeal_samples[2540]=17797;
squeal_samples[2541]=20619;
squeal_samples[2542]=23325;
squeal_samples[2543]=25907;
squeal_samples[2544]=28379;
squeal_samples[2545]=30738;
squeal_samples[2546]=32999;
squeal_samples[2547]=35154;
squeal_samples[2548]=37224;
squeal_samples[2549]=39186;
squeal_samples[2550]=41077;
squeal_samples[2551]=42869;
squeal_samples[2552]=44593;
squeal_samples[2553]=46231;
squeal_samples[2554]=47803;
squeal_samples[2555]=49301;
squeal_samples[2556]=50736;
squeal_samples[2557]=49606;
squeal_samples[2558]=44669;
squeal_samples[2559]=39998;
squeal_samples[2560]=35629;
squeal_samples[2561]=31540;
squeal_samples[2562]=27716;
squeal_samples[2563]=24139;
squeal_samples[2564]=20787;
squeal_samples[2565]=17653;
squeal_samples[2566]=14726;
squeal_samples[2567]=11986;
squeal_samples[2568]=9428;
squeal_samples[2569]=8120;
squeal_samples[2570]=10965;
squeal_samples[2571]=14079;
squeal_samples[2572]=17059;
squeal_samples[2573]=19919;
squeal_samples[2574]=22647;
squeal_samples[2575]=25261;
squeal_samples[2576]=27762;
squeal_samples[2577]=30144;
squeal_samples[2578]=32432;
squeal_samples[2579]=34610;
squeal_samples[2580]=36699;
squeal_samples[2581]=38686;
squeal_samples[2582]=40596;
squeal_samples[2583]=42416;
squeal_samples[2584]=44156;
squeal_samples[2585]=45817;
squeal_samples[2586]=47402;
squeal_samples[2587]=48921;
squeal_samples[2588]=50366;
squeal_samples[2589]=50473;
squeal_samples[2590]=45875;
squeal_samples[2591]=41124;
squeal_samples[2592]=36681;
squeal_samples[2593]=32521;
squeal_samples[2594]=28637;
squeal_samples[2595]=24999;
squeal_samples[2596]=21594;
squeal_samples[2597]=18407;
squeal_samples[2598]=15422;
squeal_samples[2599]=12644;
squeal_samples[2600]=10032;
squeal_samples[2601]=7995;
squeal_samples[2602]=10156;
squeal_samples[2603]=13301;
squeal_samples[2604]=16312;
squeal_samples[2605]=19200;
squeal_samples[2606]=21961;
squeal_samples[2607]=24605;
squeal_samples[2608]=27132;
squeal_samples[2609]=29550;
squeal_samples[2610]=31853;
squeal_samples[2611]=34062;
squeal_samples[2612]=36172;
squeal_samples[2613]=38187;
squeal_samples[2614]=40115;
squeal_samples[2615]=41951;
squeal_samples[2616]=43717;
squeal_samples[2617]=45392;
squeal_samples[2618]=47002;
squeal_samples[2619]=48529;
squeal_samples[2620]=50001;
squeal_samples[2621]=50938;
squeal_samples[2622]=47094;
squeal_samples[2623]=42269;
squeal_samples[2624]=37749;
squeal_samples[2625]=33522;
squeal_samples[2626]=29576;
squeal_samples[2627]=25870;
squeal_samples[2628]=22406;
squeal_samples[2629]=19170;
squeal_samples[2630]=16138;
squeal_samples[2631]=13308;
squeal_samples[2632]=10657;
squeal_samples[2633]=8224;
squeal_samples[2634]=9335;
squeal_samples[2635]=12515;
squeal_samples[2636]=15555;
squeal_samples[2637]=18480;
squeal_samples[2638]=21269;
squeal_samples[2639]=23942;
squeal_samples[2640]=26499;
squeal_samples[2641]=28939;
squeal_samples[2642]=31275;
squeal_samples[2643]=33507;
squeal_samples[2644]=35636;
squeal_samples[2645]=37683;
squeal_samples[2646]=39625;
squeal_samples[2647]=41491;
squeal_samples[2648]=43272;
squeal_samples[2649]=44962;
squeal_samples[2650]=46591;
squeal_samples[2651]=48142;
squeal_samples[2652]=49627;
squeal_samples[2653]=50996;
squeal_samples[2654]=48340;
squeal_samples[2655]=43437;
squeal_samples[2656]=38836;
squeal_samples[2657]=34544;
squeal_samples[2658]=30515;
squeal_samples[2659]=26760;
squeal_samples[2660]=23240;
squeal_samples[2661]=19943;
squeal_samples[2662]=16864;
squeal_samples[2663]=13986;
squeal_samples[2664]=11287;
squeal_samples[2665]=8776;
squeal_samples[2666]=8545;
squeal_samples[2667]=11721;
squeal_samples[2668]=14792;
squeal_samples[2669]=17744;
squeal_samples[2670]=20567;
squeal_samples[2671]=23271;
squeal_samples[2672]=25854;
squeal_samples[2673]=28327;
squeal_samples[2674]=30683;
squeal_samples[2675]=32949;
squeal_samples[2676]=35099;
squeal_samples[2677]=37170;
squeal_samples[2678]=39136;
squeal_samples[2679]=41020;
squeal_samples[2680]=42820;
squeal_samples[2681]=44536;
squeal_samples[2682]=46181;
squeal_samples[2683]=47748;
squeal_samples[2684]=49249;
squeal_samples[2685]=50683;
squeal_samples[2686]=49550;
squeal_samples[2687]=44619;
squeal_samples[2688]=39943;
squeal_samples[2689]=35576;
squeal_samples[2690]=31488;
squeal_samples[2691]=27663;
squeal_samples[2692]=24084;
squeal_samples[2693]=20735;
squeal_samples[2694]=17599;
squeal_samples[2695]=14673;
squeal_samples[2696]=11935;
squeal_samples[2697]=9372;
squeal_samples[2698]=8069;
squeal_samples[2699]=10910;
squeal_samples[2700]=14026;
squeal_samples[2701]=17008;
squeal_samples[2702]=19863;
squeal_samples[2703]=22597;
squeal_samples[2704]=25204;
squeal_samples[2705]=27712;
squeal_samples[2706]=30089;
squeal_samples[2707]=32379;
squeal_samples[2708]=34558;
squeal_samples[2709]=36644;
squeal_samples[2710]=38634;
squeal_samples[2711]=40542;
squeal_samples[2712]=42363;
squeal_samples[2713]=44102;
squeal_samples[2714]=45765;
squeal_samples[2715]=47348;
squeal_samples[2716]=48868;
squeal_samples[2717]=50312;
squeal_samples[2718]=50422;
squeal_samples[2719]=45819;
squeal_samples[2720]=41073;
squeal_samples[2721]=36626;
squeal_samples[2722]=32468;
squeal_samples[2723]=28585;
squeal_samples[2724]=24945;
squeal_samples[2725]=21541;
squeal_samples[2726]=18352;
squeal_samples[2727]=15370;
squeal_samples[2728]=12592;
squeal_samples[2729]=9976;
squeal_samples[2730]=7944;
squeal_samples[2731]=10101;
squeal_samples[2732]=13248;
squeal_samples[2733]=16260;
squeal_samples[2734]=19145;
squeal_samples[2735]=21909;
squeal_samples[2736]=24552;
squeal_samples[2737]=27077;
squeal_samples[2738]=29498;
squeal_samples[2739]=31799;
squeal_samples[2740]=34009;
squeal_samples[2741]=36119;
squeal_samples[2742]=38134;
squeal_samples[2743]=40060;
squeal_samples[2744]=41901;
squeal_samples[2745]=43658;
squeal_samples[2746]=45344;
squeal_samples[2747]=46945;
squeal_samples[2748]=48478;
squeal_samples[2749]=49947;
squeal_samples[2750]=50883;
squeal_samples[2751]=47042;
squeal_samples[2752]=42215;
squeal_samples[2753]=37696;
squeal_samples[2754]=33468;
squeal_samples[2755]=29524;
squeal_samples[2756]=25814;
squeal_samples[2757]=22357;
squeal_samples[2758]=19111;
squeal_samples[2759]=16089;
squeal_samples[2760]=13252;
squeal_samples[2761]=10606;
squeal_samples[2762]=8168;
squeal_samples[2763]=9285;
squeal_samples[2764]=12456;
squeal_samples[2765]=15508;
squeal_samples[2766]=18422;
squeal_samples[2767]=21218;
squeal_samples[2768]=23887;
squeal_samples[2769]=26445;
squeal_samples[2770]=28887;
squeal_samples[2771]=31222;
squeal_samples[2772]=33451;
squeal_samples[2773]=35586;
squeal_samples[2774]=37624;
squeal_samples[2775]=39578;
squeal_samples[2776]=41433;
squeal_samples[2777]=43220;
squeal_samples[2778]=44908;
squeal_samples[2779]=46537;
squeal_samples[2780]=48088;
squeal_samples[2781]=49575;
squeal_samples[2782]=50986;
squeal_samples[2783]=49091;
squeal_samples[2784]=44123;
squeal_samples[2785]=39486;
squeal_samples[2786]=35146;
squeal_samples[2787]=31075;
squeal_samples[2788]=27284;
squeal_samples[2789]=23720;
squeal_samples[2790]=20398;
squeal_samples[2791]=17281;
squeal_samples[2792]=14373;
squeal_samples[2793]=11648;
squeal_samples[2794]=9099;
squeal_samples[2795]=8293;
squeal_samples[2796]=11339;
squeal_samples[2797]=14431;
squeal_samples[2798]=17395;
squeal_samples[2799]=20232;
squeal_samples[2800]=22945;
squeal_samples[2801]=25542;
squeal_samples[2802]=28025;
squeal_samples[2803]=30396;
squeal_samples[2804]=32659;
squeal_samples[2805]=34838;
squeal_samples[2806]=36897;
squeal_samples[2807]=38886;
squeal_samples[2808]=40774;
squeal_samples[2809]=42587;
squeal_samples[2810]=44309;
squeal_samples[2811]=45964;
squeal_samples[2812]=47536;
squeal_samples[2813]=49044;
squeal_samples[2814]=50484;
squeal_samples[2815]=50581;
squeal_samples[2816]=45965;
squeal_samples[2817]=41205;
squeal_samples[2818]=36749;
squeal_samples[2819]=32580;
squeal_samples[2820]=28683;
squeal_samples[2821]=25039;
squeal_samples[2822]=21616;
squeal_samples[2823]=18430;
squeal_samples[2824]=15434;
squeal_samples[2825]=12650;
squeal_samples[2826]=10036;
squeal_samples[2827]=7992;
squeal_samples[2828]=10146;
squeal_samples[2829]=13286;
squeal_samples[2830]=16298;
squeal_samples[2831]=19179;
squeal_samples[2832]=21940;
squeal_samples[2833]=24575;
squeal_samples[2834]=27105;
squeal_samples[2835]=29515;
squeal_samples[2836]=31820;
squeal_samples[2837]=34021;
squeal_samples[2838]=36133;
squeal_samples[2839]=38149;
squeal_samples[2840]=40067;
squeal_samples[2841]=41911;
squeal_samples[2842]=43661;
squeal_samples[2843]=45345;
squeal_samples[2844]=46950;
squeal_samples[2845]=48478;
squeal_samples[2846]=49947;
squeal_samples[2847]=51135;
squeal_samples[2848]=47821;
squeal_samples[2849]=42943;
squeal_samples[2850]=38374;
squeal_samples[2851]=34107;
squeal_samples[2852]=30101;
squeal_samples[2853]=26372;
squeal_samples[2854]=22865;
squeal_samples[2855]=19591;
squeal_samples[2856]=16530;
squeal_samples[2857]=13663;
squeal_samples[2858]=10988;
squeal_samples[2859]=8479;
squeal_samples[2860]=8924;
squeal_samples[2861]=12118;
squeal_samples[2862]=15173;
squeal_samples[2863]=18105;
squeal_samples[2864]=20908;
squeal_samples[2865]=23594;
squeal_samples[2866]=26158;
squeal_samples[2867]=28616;
squeal_samples[2868]=30951;
squeal_samples[2869]=33202;
squeal_samples[2870]=35343;
squeal_samples[2871]=37390;
squeal_samples[2872]=39351;
squeal_samples[2873]=41215;
squeal_samples[2874]=43005;
squeal_samples[2875]=44713;
squeal_samples[2876]=46342;
squeal_samples[2877]=47903;
squeal_samples[2878]=49391;
squeal_samples[2879]=50812;
squeal_samples[2880]=49676;
squeal_samples[2881]=44717;
squeal_samples[2882]=40045;
squeal_samples[2883]=35658;
squeal_samples[2884]=31558;
squeal_samples[2885]=27732;
squeal_samples[2886]=24137;
squeal_samples[2887]=20781;
squeal_samples[2888]=17637;
squeal_samples[2889]=14702;
squeal_samples[2890]=11956;
squeal_samples[2891]=9386;
squeal_samples[2892]=8079;
squeal_samples[2893]=10918;
squeal_samples[2894]=14026;
squeal_samples[2895]=17009;
squeal_samples[2896]=19860;
squeal_samples[2897]=22585;
squeal_samples[2898]=25197;
squeal_samples[2899]=27693;
squeal_samples[2900]=30078;
squeal_samples[2901]=32355;
squeal_samples[2902]=34540;
squeal_samples[2903]=36616;
squeal_samples[2904]=38609;
squeal_samples[2905]=40516;
squeal_samples[2906]=42330;
squeal_samples[2907]=44068;
squeal_samples[2908]=45724;
squeal_samples[2909]=47314;
squeal_samples[2910]=48823;
squeal_samples[2911]=50272;
squeal_samples[2912]=50833;
squeal_samples[2913]=46550;
squeal_samples[2914]=41746;
squeal_samples[2915]=37254;
squeal_samples[2916]=33055;
squeal_samples[2917]=29123;
squeal_samples[2918]=25447;
squeal_samples[2919]=22001;
squeal_samples[2920]=18780;
squeal_samples[2921]=15766;
squeal_samples[2922]=12951;
squeal_samples[2923]=10317;
squeal_samples[2924]=8029;
squeal_samples[2925]=9708;
squeal_samples[2926]=12866;
squeal_samples[2927]=15895;
squeal_samples[2928]=18785;
squeal_samples[2929]=21565;
squeal_samples[2930]=24214;
squeal_samples[2931]=26761;
squeal_samples[2932]=29182;
squeal_samples[2933]=31497;
squeal_samples[2934]=33718;
squeal_samples[2935]=35836;
squeal_samples[2936]=37866;
squeal_samples[2937]=39792;
squeal_samples[2938]=41650;
squeal_samples[2939]=43408;
squeal_samples[2940]=45103;
squeal_samples[2941]=46710;
squeal_samples[2942]=48251;
squeal_samples[2943]=49725;
squeal_samples[2944]=51080;
squeal_samples[2945]=48418;
squeal_samples[2946]=43499;
squeal_samples[2947]=38891;
squeal_samples[2948]=34585;
squeal_samples[2949]=30548;
squeal_samples[2950]=26781;
squeal_samples[2951]=23249;
squeal_samples[2952]=19949;
squeal_samples[2953]=16857;
squeal_samples[2954]=13975;
squeal_samples[2955]=11270;
squeal_samples[2956]=8747;
squeal_samples[2957]=8518;
squeal_samples[2958]=11687;
squeal_samples[2959]=14761;
squeal_samples[2960]=17703;
squeal_samples[2961]=20524;
squeal_samples[2962]=23220;
squeal_samples[2963]=25807;
squeal_samples[2964]=28275;
squeal_samples[2965]=30625;
squeal_samples[2966]=32884;
squeal_samples[2967]=35039;
squeal_samples[2968]=37100;
squeal_samples[2969]=39067;
squeal_samples[2970]=40948;
squeal_samples[2971]=42747;
squeal_samples[2972]=44462;
squeal_samples[2973]=46102;
squeal_samples[2974]=47672;
squeal_samples[2975]=49168;
squeal_samples[2976]=50597;
squeal_samples[2977]=50130;
squeal_samples[2978]=45288;
squeal_samples[2979]=40569;
squeal_samples[2980]=36152;
squeal_samples[2981]=32017;
squeal_samples[2982]=28159;
squeal_samples[2983]=24532;
squeal_samples[2984]=21154;
squeal_samples[2985]=17979;
squeal_samples[2986]=15019;
squeal_samples[2987]=12250;
squeal_samples[2988]=9659;
squeal_samples[2989]=7944;
squeal_samples[2990]=10481;
squeal_samples[2991]=13605;
squeal_samples[2992]=16603;
squeal_samples[2993]=19463;
squeal_samples[2994]=22218;
squeal_samples[2995]=24834;
squeal_samples[2996]=27353;
squeal_samples[2997]=29741;
squeal_samples[2998]=32039;
squeal_samples[2999]=34222;
squeal_samples[3000]=36327;
squeal_samples[3001]=38323;
squeal_samples[3002]=40241;
squeal_samples[3003]=42072;
squeal_samples[3004]=43813;
squeal_samples[3005]=45481;
squeal_samples[3006]=47077;
squeal_samples[3007]=48599;
squeal_samples[3008]=50058;
squeal_samples[3009]=50983;
squeal_samples[3010]=47132;
squeal_samples[3011]=42291;
squeal_samples[3012]=37764;
squeal_samples[3013]=33526;
squeal_samples[3014]=29561;
squeal_samples[3015]=25852;
squeal_samples[3016]=22378;
squeal_samples[3017]=19126;
squeal_samples[3018]=16096;
squeal_samples[3019]=13249;
squeal_samples[3020]=10602;
squeal_samples[3021]=8156;
squeal_samples[3022]=9267;
squeal_samples[3023]=12435;
squeal_samples[3024]=15480;
squeal_samples[3025]=18394;
squeal_samples[3026]=21187;
squeal_samples[3027]=23851;
squeal_samples[3028]=26410;
squeal_samples[3029]=28845;
squeal_samples[3030]=31176;
squeal_samples[3031]=33404;
squeal_samples[3032]=35540;
squeal_samples[3033]=37574;
squeal_samples[3034]=39516;
squeal_samples[3035]=41381;
squeal_samples[3036]=43152;
squeal_samples[3037]=44856;
squeal_samples[3038]=46471;
squeal_samples[3039]=48026;
squeal_samples[3040]=49506;
squeal_samples[3041]=50922;
squeal_samples[3042]=49012;
squeal_samples[3043]=44061;
squeal_samples[3044]=39407;
squeal_samples[3045]=35070;
squeal_samples[3046]=30996;
squeal_samples[3047]=27204;
squeal_samples[3048]=23638;
squeal_samples[3049]=20312;
squeal_samples[3050]=17192;
squeal_samples[3051]=14282;
squeal_samples[3052]=11560;
squeal_samples[3053]=9014;
squeal_samples[3054]=8204;
squeal_samples[3055]=11249;
squeal_samples[3056]=14341;
squeal_samples[3057]=17307;
squeal_samples[3058]=20141;
squeal_samples[3059]=22857;
squeal_samples[3060]=25450;
squeal_samples[3061]=27934;
squeal_samples[3062]=30296;
squeal_samples[3063]=32571;
squeal_samples[3064]=34735;
squeal_samples[3065]=36810;
squeal_samples[3066]=38784;
squeal_samples[3067]=40680;
squeal_samples[3068]=42482;
squeal_samples[3069]=44213;
squeal_samples[3070]=45860;
squeal_samples[3071]=47437;
squeal_samples[3072]=48944;
squeal_samples[3073]=50384;
squeal_samples[3074]=50481;
squeal_samples[3075]=45865;
squeal_samples[3076]=41102;
squeal_samples[3077]=36653;
squeal_samples[3078]=32476;
squeal_samples[3079]=28587;
squeal_samples[3080]=24935;
squeal_samples[3081]=21519;
squeal_samples[3082]=18326;
squeal_samples[3083]=15339;
squeal_samples[3084]=12546;
squeal_samples[3085]=9932;
squeal_samples[3086]=7887;
squeal_samples[3087]=10045;
squeal_samples[3088]=13187;
squeal_samples[3089]=16196;
squeal_samples[3090]=19081;
squeal_samples[3091]=21838;
squeal_samples[3092]=24478;
squeal_samples[3093]=27002;
squeal_samples[3094]=29410;
squeal_samples[3095]=31721;
squeal_samples[3096]=33920;
squeal_samples[3097]=36030;
squeal_samples[3098]=38040;
squeal_samples[3099]=39970;
squeal_samples[3100]=41803;
squeal_samples[3101]=43563;
squeal_samples[3102]=45240;
squeal_samples[3103]=46844;
squeal_samples[3104]=48373;
squeal_samples[3105]=49841;
squeal_samples[3106]=51029;
squeal_samples[3107]=47724;
squeal_samples[3108]=42839;
squeal_samples[3109]=38274;
squeal_samples[3110]=33996;
squeal_samples[3111]=30000;
squeal_samples[3112]=26265;
squeal_samples[3113]=22759;
squeal_samples[3114]=19488;
squeal_samples[3115]=16421;
squeal_samples[3116]=13561;
squeal_samples[3117]=10881;
squeal_samples[3118]=8374;
squeal_samples[3119]=8820;
squeal_samples[3120]=12009;
squeal_samples[3121]=15072;
squeal_samples[3122]=17996;
squeal_samples[3123]=20806;
squeal_samples[3124]=23486;
squeal_samples[3125]=26056;
squeal_samples[3126]=28507;
squeal_samples[3127]=30849;
squeal_samples[3128]=33094;
squeal_samples[3129]=35240;
squeal_samples[3130]=37285;
squeal_samples[3131]=39243;
squeal_samples[3132]=41113;
squeal_samples[3133]=42897;
squeal_samples[3134]=44609;
squeal_samples[3135]=46236;
squeal_samples[3136]=47798;
squeal_samples[3137]=49285;
squeal_samples[3138]=50707;
squeal_samples[3139]=50227;
squeal_samples[3140]=45377;
squeal_samples[3141]=40655;
squeal_samples[3142]=36216;
squeal_samples[3143]=32083;
squeal_samples[3144]=28207;
squeal_samples[3145]=24585;
squeal_samples[3146]=21189;
squeal_samples[3147]=18011;
squeal_samples[3148]=15047;
squeal_samples[3149]=12271;
squeal_samples[3150]=9668;
squeal_samples[3151]=7952;
squeal_samples[3152]=10482;
squeal_samples[3153]=13614;
squeal_samples[3154]=16599;
squeal_samples[3155]=19467;
squeal_samples[3156]=22208;
squeal_samples[3157]=24833;
squeal_samples[3158]=27336;
squeal_samples[3159]=29731;
squeal_samples[3160]=32020;
squeal_samples[3161]=34215;
squeal_samples[3162]=36301;
squeal_samples[3163]=38307;
squeal_samples[3164]=40211;
squeal_samples[3165]=42045;
squeal_samples[3166]=43785;
squeal_samples[3167]=45454;
squeal_samples[3168]=47043;
squeal_samples[3169]=48567;
squeal_samples[3170]=50023;
squeal_samples[3171]=51207;
squeal_samples[3172]=47879;
squeal_samples[3173]=42990;
squeal_samples[3174]=38412;
squeal_samples[3175]=34131;
squeal_samples[3176]=30118;
squeal_samples[3177]=26375;
squeal_samples[3178]=22859;
squeal_samples[3179]=19579;
squeal_samples[3180]=16506;
squeal_samples[3181]=13636;
squeal_samples[3182]=10953;
squeal_samples[3183]=8441;
squeal_samples[3184]=8878;
squeal_samples[3185]=12069;
squeal_samples[3186]=15117;
squeal_samples[3187]=18049;
squeal_samples[3188]=20849;
squeal_samples[3189]=23531;
squeal_samples[3190]=26094;
squeal_samples[3191]=28548;
squeal_samples[3192]=30886;
squeal_samples[3193]=33124;
squeal_samples[3194]=35267;
squeal_samples[3195]=37312;
squeal_samples[3196]=39269;
squeal_samples[3197]=41134;
squeal_samples[3198]=42919;
squeal_samples[3199]=44628;
squeal_samples[3200]=46252;
squeal_samples[3201]=47811;
squeal_samples[3202]=49297;
squeal_samples[3203]=50718;
squeal_samples[3204]=50238;
squeal_samples[3205]=45388;
squeal_samples[3206]=40656;
squeal_samples[3207]=36223;
squeal_samples[3208]=32078;
squeal_samples[3209]=28207;
squeal_samples[3210]=24580;
squeal_samples[3211]=21183;
squeal_samples[3212]=18010;
squeal_samples[3213]=15035;
squeal_samples[3214]=12261;
squeal_samples[3215]=9661;
squeal_samples[3216]=7939;
squeal_samples[3217]=10475;
squeal_samples[3218]=13599;
squeal_samples[3219]=16587;
squeal_samples[3220]=19453;
squeal_samples[3221]=22194;
squeal_samples[3222]=24815;
squeal_samples[3223]=27326;
squeal_samples[3224]=29710;
squeal_samples[3225]=32011;
squeal_samples[3226]=34193;
squeal_samples[3227]=36293;
squeal_samples[3228]=38286;
squeal_samples[3229]=40201;
squeal_samples[3230]=42022;
squeal_samples[3231]=43770;
squeal_samples[3232]=45440;
squeal_samples[3233]=47027;
squeal_samples[3234]=48553;
squeal_samples[3235]=50003;
squeal_samples[3236]=51184;
squeal_samples[3237]=47863;
squeal_samples[3238]=42963;
squeal_samples[3239]=38394;
squeal_samples[3240]=34103;
squeal_samples[3241]=30098;
squeal_samples[3242]=26350;
squeal_samples[3243]=22842;
squeal_samples[3244]=19556;
squeal_samples[3245]=16488;
squeal_samples[3246]=13608;
squeal_samples[3247]=10929;
squeal_samples[3248]=8419;
squeal_samples[3249]=8855;
squeal_samples[3250]=12039;
squeal_samples[3251]=15101;
squeal_samples[3252]=18025;
squeal_samples[3253]=20826;
squeal_samples[3254]=23504;
squeal_samples[3255]=26068;
squeal_samples[3256]=28523;
squeal_samples[3257]=30859;
squeal_samples[3258]=33105;
squeal_samples[3259]=35240;
squeal_samples[3260]=37287;
squeal_samples[3261]=39243;
squeal_samples[3262]=41107;
squeal_samples[3263]=42896;
squeal_samples[3264]=44600;
squeal_samples[3265]=46228;
squeal_samples[3266]=47783;
squeal_samples[3267]=49272;
squeal_samples[3268]=50694;
squeal_samples[3269]=50211;
squeal_samples[3270]=45363;
squeal_samples[3271]=40629;
squeal_samples[3272]=36204;
squeal_samples[3273]=32052;
squeal_samples[3274]=28182;
squeal_samples[3275]=24552;
squeal_samples[3276]=21160;
squeal_samples[3277]=17982;
squeal_samples[3278]=15010;
squeal_samples[3279]=12236;
squeal_samples[3280]=9634;
squeal_samples[3281]=7915;
squeal_samples[3282]=10448;
squeal_samples[3283]=13578;
squeal_samples[3284]=16564;
squeal_samples[3285]=19425;
squeal_samples[3286]=22170;
squeal_samples[3287]=24789;
squeal_samples[3288]=27299;
squeal_samples[3289]=29686;
squeal_samples[3290]=31984;
squeal_samples[3291]=34168;
squeal_samples[3292]=36268;
squeal_samples[3293]=38260;
squeal_samples[3294]=40175;
squeal_samples[3295]=41995;
squeal_samples[3296]=43747;
squeal_samples[3297]=45412;
squeal_samples[3298]=47002;
squeal_samples[3299]=48529;
squeal_samples[3300]=49973;
squeal_samples[3301]=51165;
squeal_samples[3302]=47830;
squeal_samples[3303]=42945;
squeal_samples[3304]=38366;
squeal_samples[3305]=34083;
squeal_samples[3306]=30070;
squeal_samples[3307]=26325;
squeal_samples[3308]=22817;
squeal_samples[3309]=19529;
squeal_samples[3310]=16463;
squeal_samples[3311]=13583;
squeal_samples[3312]=10902;
squeal_samples[3313]=8395;
squeal_samples[3314]=8827;
squeal_samples[3315]=12017;
squeal_samples[3316]=15071;
squeal_samples[3317]=18004;
squeal_samples[3318]=20796;
squeal_samples[3319]=23482;
squeal_samples[3320]=26041;
squeal_samples[3321]=28496;
squeal_samples[3322]=30836;
squeal_samples[3323]=33077;
squeal_samples[3324]=35216;
squeal_samples[3325]=37262;
squeal_samples[3326]=39215;
squeal_samples[3327]=41083;
squeal_samples[3328]=42871;
squeal_samples[3329]=44571;
squeal_samples[3330]=46207;
squeal_samples[3331]=47754;
squeal_samples[3332]=49248;
squeal_samples[3333]=50668;
squeal_samples[3334]=50184;
squeal_samples[3335]=45339;
squeal_samples[3336]=40603;
squeal_samples[3337]=36177;
squeal_samples[3338]=32028;
squeal_samples[3339]=28155;
squeal_samples[3340]=24527;
squeal_samples[3341]=21135;
squeal_samples[3342]=17955;
squeal_samples[3343]=14987;
squeal_samples[3344]=12207;
squeal_samples[3345]=9612;
squeal_samples[3346]=7886;
squeal_samples[3347]=10425;
squeal_samples[3348]=13552;
squeal_samples[3349]=16537;
squeal_samples[3350]=19401;
squeal_samples[3351]=22143;
squeal_samples[3352]=24764;
squeal_samples[3353]=27274;
squeal_samples[3354]=29660;
squeal_samples[3355]=31958;
squeal_samples[3356]=34144;
squeal_samples[3357]=36238;
squeal_samples[3358]=38240;
squeal_samples[3359]=40145;
squeal_samples[3360]=41973;
squeal_samples[3361]=43720;
squeal_samples[3362]=45385;
squeal_samples[3363]=46980;
squeal_samples[3364]=48499;
squeal_samples[3365]=49952;
squeal_samples[3366]=51135;
squeal_samples[3367]=47809;
squeal_samples[3368]=42915;
squeal_samples[3369]=38345;
squeal_samples[3370]=34054;
squeal_samples[3371]=30046;
squeal_samples[3372]=26300;
squeal_samples[3373]=22788;
squeal_samples[3374]=19509;
squeal_samples[3375]=16431;
squeal_samples[3376]=13563;
squeal_samples[3377]=10875;
squeal_samples[3378]=8367;
squeal_samples[3379]=8806;
squeal_samples[3380]=11986;
squeal_samples[3381]=15051;
squeal_samples[3382]=17974;
squeal_samples[3383]=20774;
squeal_samples[3384]=23452;
squeal_samples[3385]=26020;
squeal_samples[3386]=28468;
squeal_samples[3387]=30812;
squeal_samples[3388]=33051;
squeal_samples[3389]=35189;
squeal_samples[3390]=37238;
squeal_samples[3391]=39189;
squeal_samples[3392]=41059;
squeal_samples[3393]=42843;
squeal_samples[3394]=44548;
squeal_samples[3395]=46179;
squeal_samples[3396]=47731;
squeal_samples[3397]=49222;
squeal_samples[3398]=50641;
squeal_samples[3399]=50160;
squeal_samples[3400]=45312;
squeal_samples[3401]=40579;
squeal_samples[3402]=36151;
squeal_samples[3403]=32002;
squeal_samples[3404]=28130;
squeal_samples[3405]=24502;
squeal_samples[3406]=21108;
squeal_samples[3407]=17931;
squeal_samples[3408]=14959;
squeal_samples[3409]=12184;
squeal_samples[3410]=9585;
squeal_samples[3411]=7861;
squeal_samples[3412]=10399;
squeal_samples[3413]=13527;
squeal_samples[3414]=16511;
squeal_samples[3415]=19376;
squeal_samples[3416]=22117;
squeal_samples[3417]=24739;
squeal_samples[3418]=27248;
squeal_samples[3419]=29635;
squeal_samples[3420]=31932;
squeal_samples[3421]=34118;
squeal_samples[3422]=36216;
squeal_samples[3423]=38210;
squeal_samples[3424]=40123;
squeal_samples[3425]=41945;
squeal_samples[3426]=43695;
squeal_samples[3427]=45361;
squeal_samples[3428]=46954;
squeal_samples[3429]=48473;
squeal_samples[3430]=49926;
squeal_samples[3431]=51112;
squeal_samples[3432]=47779;
squeal_samples[3433]=42895;
squeal_samples[3434]=38315;
squeal_samples[3435]=34031;
squeal_samples[3436]=30020;
squeal_samples[3437]=26274;
squeal_samples[3438]=22764;
squeal_samples[3439]=19481;
squeal_samples[3440]=16409;
squeal_samples[3441]=13534;
squeal_samples[3442]=10851;
squeal_samples[3443]=8343;
squeal_samples[3444]=8777;
squeal_samples[3445]=11964;
squeal_samples[3446]=15022;
squeal_samples[3447]=17952;
squeal_samples[3448]=20745;
squeal_samples[3449]=23431;
squeal_samples[3450]=25990;
squeal_samples[3451]=28445;
squeal_samples[3452]=30785;
squeal_samples[3453]=33025;
squeal_samples[3454]=35167;
squeal_samples[3455]=37208;
squeal_samples[3456]=39168;
squeal_samples[3457]=41029;
squeal_samples[3458]=42821;
squeal_samples[3459]=44521;
squeal_samples[3460]=46154;
squeal_samples[3461]=47705;
squeal_samples[3462]=49197;
squeal_samples[3463]=50615;
squeal_samples[3464]=50136;
squeal_samples[3465]=45285;
squeal_samples[3466]=40554;
squeal_samples[3467]=36126;
squeal_samples[3468]=31976;
squeal_samples[3469]=28105;
squeal_samples[3470]=24476;
squeal_samples[3471]=21082;
squeal_samples[3472]=17908;
squeal_samples[3473]=14931;
squeal_samples[3474]=12161;
squeal_samples[3475]=9558;
squeal_samples[3476]=7835;
squeal_samples[3477]=10375;
squeal_samples[3478]=13500;
squeal_samples[3479]=16487;
squeal_samples[3480]=19350;
squeal_samples[3481]=22091;
squeal_samples[3482]=24713;
squeal_samples[3483]=27224;
squeal_samples[3484]=29608;
squeal_samples[3485]=31907;
squeal_samples[3486]=34093;
squeal_samples[3487]=36189;
squeal_samples[3488]=38185;
squeal_samples[3489]=40099;
squeal_samples[3490]=41917;
squeal_samples[3491]=43671;
squeal_samples[3492]=45333;
squeal_samples[3493]=46930;
squeal_samples[3494]=48446;
squeal_samples[3495]=49903;
squeal_samples[3496]=51238;
squeal_samples[3497]=48557;
squeal_samples[3498]=43610;
squeal_samples[3499]=38986;
squeal_samples[3500]=34658;
squeal_samples[3501]=30605;
squeal_samples[3502]=26822;
squeal_samples[3503]=23267;
squeal_samples[3504]=19953;
squeal_samples[3505]=16846;
squeal_samples[3506]=13953;
squeal_samples[3507]=11229;
squeal_samples[3508]=8701;
squeal_samples[3509]=8461;
squeal_samples[3510]=11619;
squeal_samples[3511]=14686;
squeal_samples[3512]=17628;
squeal_samples[3513]=20437;
squeal_samples[3514]=23133;
squeal_samples[3515]=25710;
squeal_samples[3516]=28175;
squeal_samples[3517]=30521;
squeal_samples[3518]=32772;
squeal_samples[3519]=34921;
squeal_samples[3520]=36980;
squeal_samples[3521]=38943;
squeal_samples[3522]=40822;
squeal_samples[3523]=42614;
squeal_samples[3524]=44323;
squeal_samples[3525]=45963;
squeal_samples[3526]=47524;
squeal_samples[3527]=49016;
squeal_samples[3528]=50449;
squeal_samples[3529]=50990;
squeal_samples[3530]=46677;
squeal_samples[3531]=41854;
squeal_samples[3532]=37339;
squeal_samples[3533]=33112;
squeal_samples[3534]=29165;
squeal_samples[3535]=25467;
squeal_samples[3536]=22006;
squeal_samples[3537]=18772;
squeal_samples[3538]=15739;
squeal_samples[3539]=12907;
squeal_samples[3540]=10267;
squeal_samples[3541]=7962;
squeal_samples[3542]=9636;
squeal_samples[3543]=12780;
squeal_samples[3544]=15807;
squeal_samples[3545]=18692;
squeal_samples[3546]=21465;
squeal_samples[3547]=24111;
squeal_samples[3548]=26643;
squeal_samples[3549]=29064;
squeal_samples[3550]=31374;
squeal_samples[3551]=33587;
squeal_samples[3552]=35699;
squeal_samples[3553]=37722;
squeal_samples[3554]=39653;
squeal_samples[3555]=41497;
squeal_samples[3556]=43260;
squeal_samples[3557]=44937;
squeal_samples[3558]=46552;
squeal_samples[3559]=48083;
squeal_samples[3560]=49556;
squeal_samples[3561]=50956;
squeal_samples[3562]=49800;
squeal_samples[3563]=44821;
squeal_samples[3564]=40119;
squeal_samples[3565]=35713;
squeal_samples[3566]=31590;
squeal_samples[3567]=27740;
squeal_samples[3568]=24134;
squeal_samples[3569]=20756;
squeal_samples[3570]=17601;
squeal_samples[3571]=14646;
squeal_samples[3572]=11886;
squeal_samples[3573]=9303;
squeal_samples[3574]=7986;
squeal_samples[3575]=10821;
squeal_samples[3576]=13923;
squeal_samples[3577]=16894;
squeal_samples[3578]=19735;
squeal_samples[3579]=22460;
squeal_samples[3580]=25059;
squeal_samples[3581]=27557;
squeal_samples[3582]=29924;
squeal_samples[3583]=32210;
squeal_samples[3584]=34376;
squeal_samples[3585]=36463;
squeal_samples[3586]=38444;
squeal_samples[3587]=40342;
squeal_samples[3588]=42152;
squeal_samples[3589]=43885;
squeal_samples[3590]=45544;
squeal_samples[3591]=47119;
squeal_samples[3592]=48636;
squeal_samples[3593]=50077;
squeal_samples[3594]=51253;
squeal_samples[3595]=47914;
squeal_samples[3596]=43006;
squeal_samples[3597]=38422;
squeal_samples[3598]=34124;
squeal_samples[3599]=30106;
squeal_samples[3600]=26349;
squeal_samples[3601]=22828;
squeal_samples[3602]=19538;
squeal_samples[3603]=16458;
squeal_samples[3604]=13580;
squeal_samples[3605]=10883;
squeal_samples[3606]=8373;
squeal_samples[3607]=8799;
squeal_samples[3608]=11988;
squeal_samples[3609]=15040;
squeal_samples[3610]=17961;
squeal_samples[3611]=20761;
squeal_samples[3612]=23434;
squeal_samples[3613]=25999;
squeal_samples[3614]=28446;
squeal_samples[3615]=30779;
squeal_samples[3616]=33024;
squeal_samples[3617]=35153;
squeal_samples[3618]=37203;
squeal_samples[3619]=39154;
squeal_samples[3620]=41016;
squeal_samples[3621]=42805;
squeal_samples[3622]=44502;
squeal_samples[3623]=46132;
squeal_samples[3624]=47686;
squeal_samples[3625]=49167;
squeal_samples[3626]=50592;
squeal_samples[3627]=50662;
squeal_samples[3628]=46028;
squeal_samples[3629]=41238;
squeal_samples[3630]=36761;
squeal_samples[3631]=32578;
squeal_samples[3632]=28656;
squeal_samples[3633]=24992;
squeal_samples[3634]=21554;
squeal_samples[3635]=18347;
squeal_samples[3636]=15343;
squeal_samples[3637]=12534;
squeal_samples[3638]=9909;
squeal_samples[3639]=7852;
squeal_samples[3640]=10002;
squeal_samples[3641]=13129;
squeal_samples[3642]=16139;
squeal_samples[3643]=19011;
squeal_samples[3644]=21769;
squeal_samples[3645]=24399;
squeal_samples[3646]=26914;
squeal_samples[3647]=29324;
squeal_samples[3648]=31620;
squeal_samples[3649]=33817;
squeal_samples[3650]=35925;
squeal_samples[3651]=37930;
squeal_samples[3652]=39852;
squeal_samples[3653]=41679;
squeal_samples[3654]=43439;
squeal_samples[3655]=45108;
squeal_samples[3656]=46709;
squeal_samples[3657]=48242;
squeal_samples[3658]=49691;
squeal_samples[3659]=51099;
squeal_samples[3660]=49162;
squeal_samples[3661]=44186;
squeal_samples[3662]=39511;
squeal_samples[3663]=35152;
squeal_samples[3664]=31054;
squeal_samples[3665]=27243;
squeal_samples[3666]=23659;
squeal_samples[3667]=20318;
squeal_samples[3668]=17182;
squeal_samples[3669]=14254;
squeal_samples[3670]=11516;
squeal_samples[3671]=8957;
squeal_samples[3672]=8136;
squeal_samples[3673]=11181;
squeal_samples[3674]=14259;
squeal_samples[3675]=17214;
squeal_samples[3676]=20046;
squeal_samples[3677]=22751;
squeal_samples[3678]=25343;
squeal_samples[3679]=27820;
squeal_samples[3680]=30178;
squeal_samples[3681]=32444;
squeal_samples[3682]=34608;
squeal_samples[3683]=36671;
squeal_samples[3684]=38647;
squeal_samples[3685]=40535;
squeal_samples[3686]=42338;
squeal_samples[3687]=44060;
squeal_samples[3688]=45704;
squeal_samples[3689]=47280;
squeal_samples[3690]=48779;
squeal_samples[3691]=50216;
squeal_samples[3692]=51126;
squeal_samples[3693]=47248;
squeal_samples[3694]=42378;
squeal_samples[3695]=37833;
squeal_samples[3696]=33567;
squeal_samples[3697]=29587;
squeal_samples[3698]=25858;
squeal_samples[3699]=22367;
squeal_samples[3700]=19104;
squeal_samples[3701]=16049;
squeal_samples[3702]=13196;
squeal_samples[3703]=10523;
squeal_samples[3704]=8073;
squeal_samples[3705]=9171;
squeal_samples[3706]=12333;
squeal_samples[3707]=15373;
squeal_samples[3708]=18276;
squeal_samples[3709]=21063;
squeal_samples[3710]=23725;
squeal_samples[3711]=26267;
squeal_samples[3712]=28709;
squeal_samples[3713]=31027;
squeal_samples[3714]=33257;
squeal_samples[3715]=35378;
squeal_samples[3716]=37411;
squeal_samples[3717]=39352;
squeal_samples[3718]=41206;
squeal_samples[3719]=42982;
squeal_samples[3720]=44672;
squeal_samples[3721]=46288;
squeal_samples[3722]=47838;
squeal_samples[3723]=49311;
squeal_samples[3724]=50724;
squeal_samples[3725]=50237;
squeal_samples[3726]=45366;
squeal_samples[3727]=40626;
squeal_samples[3728]=36187;
squeal_samples[3729]=32030;
squeal_samples[3730]=28152;
squeal_samples[3731]=24507;
squeal_samples[3732]=21109;
squeal_samples[3733]=17919;
squeal_samples[3734]=14944;
squeal_samples[3735]=12157;
squeal_samples[3736]=9557;
squeal_samples[3737]=7824;
squeal_samples[3738]=10360;
squeal_samples[3739]=13479;
squeal_samples[3740]=16467;
squeal_samples[3741]=19323;
squeal_samples[3742]=22061;
squeal_samples[3743]=24681;
squeal_samples[3744]=27187;
squeal_samples[3745]=29571;
squeal_samples[3746]=31865;
squeal_samples[3747]=34052;
squeal_samples[3748]=36138;
squeal_samples[3749]=38142;
squeal_samples[3750]=40040;
squeal_samples[3751]=41870;
squeal_samples[3752]=43608;
squeal_samples[3753]=45279;
squeal_samples[3754]=46861;
squeal_samples[3755]=48386;
squeal_samples[3756]=49836;
squeal_samples[3757]=51176;
squeal_samples[3758]=48489;
squeal_samples[3759]=43537;
squeal_samples[3760]=38916;
squeal_samples[3761]=34579;
squeal_samples[3762]=30533;
squeal_samples[3763]=26740;
squeal_samples[3764]=23194;
squeal_samples[3765]=19871;
squeal_samples[3766]=16769;
squeal_samples[3767]=13864;
squeal_samples[3768]=11151;
squeal_samples[3769]=8614;
squeal_samples[3770]=8376;
squeal_samples[3771]=11533;
squeal_samples[3772]=14603;
squeal_samples[3773]=17537;
squeal_samples[3774]=20358;
squeal_samples[3775]=23041;
squeal_samples[3776]=25624;
squeal_samples[3777]=28082;
squeal_samples[3778]=30429;
squeal_samples[3779]=32682;
squeal_samples[3780]=34830;
squeal_samples[3781]=36888;
squeal_samples[3782]=38854;
squeal_samples[3783]=40724;
squeal_samples[3784]=42518;
squeal_samples[3785]=44231;
squeal_samples[3786]=45869;
squeal_samples[3787]=47430;
squeal_samples[3788]=48928;
squeal_samples[3789]=50350;
squeal_samples[3790]=50894;
squeal_samples[3791]=46582;
squeal_samples[3792]=41757;
squeal_samples[3793]=37242;
squeal_samples[3794]=33016;
squeal_samples[3795]=29069;
squeal_samples[3796]=25370;
squeal_samples[3797]=21911;
squeal_samples[3798]=18673;
squeal_samples[3799]=15644;
squeal_samples[3800]=12812;
squeal_samples[3801]=10167;
squeal_samples[3802]=7866;
squeal_samples[3803]=9532;
squeal_samples[3804]=12690;
squeal_samples[3805]=15700;
squeal_samples[3806]=18599;
squeal_samples[3807]=21361;
squeal_samples[3808]=24010;
squeal_samples[3809]=26548;
squeal_samples[3810]=28964;
squeal_samples[3811]=31276;
squeal_samples[3812]=33486;
squeal_samples[3813]=35602;
squeal_samples[3814]=37617;
squeal_samples[3815]=39552;
squeal_samples[3816]=41395;
squeal_samples[3817]=43158;
squeal_samples[3818]=44836;
squeal_samples[3819]=46447;
squeal_samples[3820]=47983;
squeal_samples[3821]=49453;
squeal_samples[3822]=50855;
squeal_samples[3823]=50359;
squeal_samples[3824]=45480;
squeal_samples[3825]=40729;
squeal_samples[3826]=36278;
squeal_samples[3827]=32120;
squeal_samples[3828]=28223;
squeal_samples[3829]=24581;
squeal_samples[3830]=21170;
squeal_samples[3831]=17976;
squeal_samples[3832]=14996;
squeal_samples[3833]=12201;
squeal_samples[3834]=9599;
squeal_samples[3835]=7857;
squeal_samples[3836]=10392;
squeal_samples[3837]=13506;
squeal_samples[3838]=16487;
squeal_samples[3839]=19351;
squeal_samples[3840]=22081;
squeal_samples[3841]=24698;
squeal_samples[3842]=27202;
squeal_samples[3843]=29588;
squeal_samples[3844]=31875;
squeal_samples[3845]=34056;
squeal_samples[3846]=36145;
squeal_samples[3847]=38144;
squeal_samples[3848]=40049;
squeal_samples[3849]=41871;
squeal_samples[3850]=43611;
squeal_samples[3851]=45270;
squeal_samples[3852]=46863;
squeal_samples[3853]=48380;
squeal_samples[3854]=49828;
squeal_samples[3855]=51168;
squeal_samples[3856]=48473;
squeal_samples[3857]=43532;
squeal_samples[3858]=38898;
squeal_samples[3859]=34568;
squeal_samples[3860]=30513;
squeal_samples[3861]=26724;
squeal_samples[3862]=23172;
squeal_samples[3863]=19855;
squeal_samples[3864]=16746;
squeal_samples[3865]=13842;
squeal_samples[3866]=11124;
squeal_samples[3867]=8585;
squeal_samples[3868]=8350;
squeal_samples[3869]=11507;
squeal_samples[3870]=14570;
squeal_samples[3871]=17517;
squeal_samples[3872]=20322;
squeal_samples[3873]=23022;
squeal_samples[3874]=25590;
squeal_samples[3875]=28053;
squeal_samples[3876]=30399;
squeal_samples[3877]=32656;
squeal_samples[3878]=34802;
squeal_samples[3879]=36856;
squeal_samples[3880]=38819;
squeal_samples[3881]=40698;
squeal_samples[3882]=42489;
squeal_samples[3883]=44200;
squeal_samples[3884]=45833;
squeal_samples[3885]=47399;
squeal_samples[3886]=48893;
squeal_samples[3887]=50317;
squeal_samples[3888]=51219;
squeal_samples[3889]=47331;
squeal_samples[3890]=42458;
squeal_samples[3891]=37892;
squeal_samples[3892]=33625;
squeal_samples[3893]=29626;
squeal_samples[3894]=25896;
squeal_samples[3895]=22401;
squeal_samples[3896]=19127;
squeal_samples[3897]=16068;
squeal_samples[3898]=13202;
squeal_samples[3899]=10531;
squeal_samples[3900]=8070;
squeal_samples[3901]=9166;
squeal_samples[3902]=12327;
squeal_samples[3903]=15365;
squeal_samples[3904]=18267;
squeal_samples[3905]=21043;
squeal_samples[3906]=23710;
squeal_samples[3907]=26249;
squeal_samples[3908]=28686;
squeal_samples[3909]=31001;
squeal_samples[3910]=33227;
squeal_samples[3911]=35350;
squeal_samples[3912]=37378;
squeal_samples[3913]=39319;
squeal_samples[3914]=41171;
squeal_samples[3915]=42945;
squeal_samples[3916]=44631;
squeal_samples[3917]=46249;
squeal_samples[3918]=47795;
squeal_samples[3919]=49264;
squeal_samples[3920]=50682;
squeal_samples[3921]=50744;
squeal_samples[3922]=46088;
squeal_samples[3923]=41300;
squeal_samples[3924]=36803;
squeal_samples[3925]=32608;
squeal_samples[3926]=28679;
squeal_samples[3927]=25004;
squeal_samples[3928]=21566;
squeal_samples[3929]=18345;
squeal_samples[3930]=15338;
squeal_samples[3931]=12520;
squeal_samples[3932]=9887;
squeal_samples[3933]=7825;
squeal_samples[3934]=9966;
squeal_samples[3935]=13099;
squeal_samples[3936]=16096;
squeal_samples[3937]=18969;
squeal_samples[3938]=21723;
squeal_samples[3939]=24351;
squeal_samples[3940]=26862;
squeal_samples[3941]=29264;
squeal_samples[3942]=31564;
squeal_samples[3943]=33762;
squeal_samples[3944]=35865;
squeal_samples[3945]=37863;
squeal_samples[3946]=39784;
squeal_samples[3947]=41615;
squeal_samples[3948]=43365;
squeal_samples[3949]=45039;
squeal_samples[3950]=46630;
squeal_samples[3951]=48164;
squeal_samples[3952]=49615;
squeal_samples[3953]=51013;
squeal_samples[3954]=49839;
squeal_samples[3955]=44853;
squeal_samples[3956]=40141;
squeal_samples[3957]=35718;
squeal_samples[3958]=31594;
squeal_samples[3959]=27724;
squeal_samples[3960]=24112;
squeal_samples[3961]=20729;
squeal_samples[3962]=17559;
squeal_samples[3963]=14602;
squeal_samples[3964]=11837;
squeal_samples[3965]=9245;
squeal_samples[3966]=7923;
squeal_samples[3967]=10752;
squeal_samples[3968]=13851;
squeal_samples[3969]=16817;
squeal_samples[3970]=19658;
squeal_samples[3971]=22376;
squeal_samples[3972]=24980;
squeal_samples[3973]=27462;
squeal_samples[3974]=29837;
squeal_samples[3975]=32111;
squeal_samples[3976]=34282;
squeal_samples[3977]=36358;
squeal_samples[3978]=38345;
squeal_samples[3979]=40232;
squeal_samples[3980]=42051;
squeal_samples[3981]=43781;
squeal_samples[3982]=45429;
squeal_samples[3983]=47015;
squeal_samples[3984]=48515;
squeal_samples[3985]=49965;
squeal_samples[3986]=51287;
squeal_samples[3987]=48592;
squeal_samples[3988]=43631;
squeal_samples[3989]=38988;
squeal_samples[3990]=34652;
squeal_samples[3991]=30588;
squeal_samples[3992]=26790;
squeal_samples[3993]=23237;
squeal_samples[3994]=19903;
squeal_samples[3995]=16795;
squeal_samples[3996]=13882;
squeal_samples[3997]=11160;
squeal_samples[3998]=8614;
squeal_samples[3999]=8376;
squeal_samples[4000]=11522;
squeal_samples[4001]=14589;
squeal_samples[4002]=17526;
squeal_samples[4003]=20334;
squeal_samples[4004]=23027;
squeal_samples[4005]=25600;
squeal_samples[4006]=28060;
squeal_samples[4007]=30404;
squeal_samples[4008]=32651;
squeal_samples[4009]=34801;
squeal_samples[4010]=36852;
squeal_samples[4011]=38812;
squeal_samples[4012]=40685;
squeal_samples[4013]=42475;
squeal_samples[4014]=44186;
squeal_samples[4015]=45820;
squeal_samples[4016]=47380;
squeal_samples[4017]=48873;
squeal_samples[4018]=50302;
squeal_samples[4019]=51196;
squeal_samples[4020]=47310;
squeal_samples[4021]=42429;
squeal_samples[4022]=37873;
squeal_samples[4023]=33592;
squeal_samples[4024]=29599;
squeal_samples[4025]=25865;
squeal_samples[4026]=22370;
squeal_samples[4027]=19094;
squeal_samples[4028]=16032;
squeal_samples[4029]=13168;
squeal_samples[4030]=10494;
squeal_samples[4031]=8037;
squeal_samples[4032]=9128;
squeal_samples[4033]=12294;
squeal_samples[4034]=15325;
squeal_samples[4035]=18224;
squeal_samples[4036]=21006;
squeal_samples[4037]=23665;
squeal_samples[4038]=26212;
squeal_samples[4039]=28644;
squeal_samples[4040]=30960;
squeal_samples[4041]=33183;
squeal_samples[4042]=35307;
squeal_samples[4043]=37340;
squeal_samples[4044]=39277;
squeal_samples[4045]=41126;
squeal_samples[4046]=42899;
squeal_samples[4047]=44588;
squeal_samples[4048]=46207;
squeal_samples[4049]=47746;
squeal_samples[4050]=49220;
squeal_samples[4051]=50636;
squeal_samples[4052]=50695;
squeal_samples[4053]=46047;
squeal_samples[4054]=41244;
squeal_samples[4055]=36761;
squeal_samples[4056]=32559;
squeal_samples[4057]=28636;
squeal_samples[4058]=24955;
squeal_samples[4059]=21518;
squeal_samples[4060]=18290;
squeal_samples[4061]=15290;
squeal_samples[4062]=12465;
squeal_samples[4063]=9845;
squeal_samples[4064]=7770;
squeal_samples[4065]=9917;
squeal_samples[4066]=13046;
squeal_samples[4067]=16051;
squeal_samples[4068]=18923;
squeal_samples[4069]=21671;
squeal_samples[4070]=24300;
squeal_samples[4071]=26816;
squeal_samples[4072]=29218;
squeal_samples[4073]=31513;
squeal_samples[4074]=33710;
squeal_samples[4075]=35813;
squeal_samples[4076]=37814;
squeal_samples[4077]=39735;
squeal_samples[4078]=41566;
squeal_samples[4079]=43313;
squeal_samples[4080]=44985;
squeal_samples[4081]=46583;
squeal_samples[4082]=48109;
squeal_samples[4083]=49566;
squeal_samples[4084]=50966;
squeal_samples[4085]=49792;
squeal_samples[4086]=44804;
squeal_samples[4087]=40086;
squeal_samples[4088]=35673;
squeal_samples[4089]=31534;
squeal_samples[4090]=27680;
squeal_samples[4091]=24056;
squeal_samples[4092]=20678;
squeal_samples[4093]=17511;
squeal_samples[4094]=14547;
squeal_samples[4095]=11786;
squeal_samples[4096]=9195;
squeal_samples[4097]=7875;
squeal_samples[4098]=10702;
squeal_samples[4099]=13800;
squeal_samples[4100]=16764;
squeal_samples[4101]=19608;
squeal_samples[4102]=22324;
squeal_samples[4103]=24928;
squeal_samples[4104]=27411;
squeal_samples[4105]=29787;
squeal_samples[4106]=32058;
squeal_samples[4107]=34230;
squeal_samples[4108]=36310;
squeal_samples[4109]=38288;
squeal_samples[4110]=40186;
squeal_samples[4111]=41997;
squeal_samples[4112]=43729;
squeal_samples[4113]=45380;
squeal_samples[4114]=46961;
squeal_samples[4115]=48465;
squeal_samples[4116]=49913;
squeal_samples[4117]=51236;
squeal_samples[4118]=48540;
squeal_samples[4119]=43580;
squeal_samples[4120]=38936;
squeal_samples[4121]=34602;
squeal_samples[4122]=30534;
squeal_samples[4123]=26740;
squeal_samples[4124]=23185;
squeal_samples[4125]=19852;
squeal_samples[4126]=16743;
squeal_samples[4127]=13831;
squeal_samples[4128]=11106;
squeal_samples[4129]=8566;
squeal_samples[4130]=8322;
squeal_samples[4131]=11472;
squeal_samples[4132]=14542;
squeal_samples[4133]=17474;
squeal_samples[4134]=20289;
squeal_samples[4135]=22975;
squeal_samples[4136]=25549;
squeal_samples[4137]=28008;
squeal_samples[4138]=30352;
squeal_samples[4139]=32600;
squeal_samples[4140]=34750;
squeal_samples[4141]=36799;
squeal_samples[4142]=38763;
squeal_samples[4143]=40630;
squeal_samples[4144]=42426;
squeal_samples[4145]=44134;
squeal_samples[4146]=45768;
squeal_samples[4147]=47330;
squeal_samples[4148]=48820;
squeal_samples[4149]=50250;
squeal_samples[4150]=51146;
squeal_samples[4151]=47256;
squeal_samples[4152]=42382;
squeal_samples[4153]=37817;
squeal_samples[4154]=33543;
squeal_samples[4155]=29546;
squeal_samples[4156]=25813;
squeal_samples[4157]=22319;
squeal_samples[4158]=19044;
squeal_samples[4159]=15978;
squeal_samples[4160]=13118;
squeal_samples[4161]=10441;
squeal_samples[4162]=7986;
squeal_samples[4163]=9077;
squeal_samples[4164]=12242;
squeal_samples[4165]=15273;
squeal_samples[4166]=18172;
squeal_samples[4167]=20956;
squeal_samples[4168]=23611;
squeal_samples[4169]=26162;
squeal_samples[4170]=28591;
squeal_samples[4171]=30910;
squeal_samples[4172]=33129;
squeal_samples[4173]=35258;
squeal_samples[4174]=37285;
squeal_samples[4175]=39226;
squeal_samples[4176]=41075;
squeal_samples[4177]=42846;
squeal_samples[4178]=44539;
squeal_samples[4179]=46153;
squeal_samples[4180]=47693;
squeal_samples[4181]=49169;
squeal_samples[4182]=50582;
squeal_samples[4183]=51108;
squeal_samples[4184]=46770;
squeal_samples[4185]=41921;
squeal_samples[4186]=37387;
squeal_samples[4187]=33143;
squeal_samples[4188]=29175;
squeal_samples[4189]=25459;
squeal_samples[4190]=21985;
squeal_samples[4191]=18730;
squeal_samples[4192]=15691;
squeal_samples[4193]=12846;
squeal_samples[4194]=10186;
squeal_samples[4195]=7873;
squeal_samples[4196]=9538;
squeal_samples[4197]=12679;
squeal_samples[4198]=15696;
squeal_samples[4199]=18575;
squeal_samples[4200]=21345;
squeal_samples[4201]=23980;
squeal_samples[4202]=26511;
squeal_samples[4203]=28927;
squeal_samples[4204]=31226;
squeal_samples[4205]=33439;
squeal_samples[4206]=35545;
squeal_samples[4207]=37565;
squeal_samples[4208]=39486;
squeal_samples[4209]=41330;
squeal_samples[4210]=43088;
squeal_samples[4211]=44764;
squeal_samples[4212]=46374;
squeal_samples[4213]=47904;
squeal_samples[4214]=49368;
squeal_samples[4215]=50771;
squeal_samples[4216]=50264;
squeal_samples[4217]=45387;
squeal_samples[4218]=40632;
squeal_samples[4219]=36179;
squeal_samples[4220]=32011;
squeal_samples[4221]=28120;
squeal_samples[4222]=24470;
squeal_samples[4223]=21052;
squeal_samples[4224]=17861;
squeal_samples[4225]=14870;
squeal_samples[4226]=12083;
squeal_samples[4227]=9470;
squeal_samples[4228]=7734;
squeal_samples[4229]=10267;
squeal_samples[4230]=13373;
squeal_samples[4231]=16367;
squeal_samples[4232]=19212;
squeal_samples[4233]=21957;
squeal_samples[4234]=24563;
squeal_samples[4235]=27069;
squeal_samples[4236]=29450;
squeal_samples[4237]=31737;
squeal_samples[4238]=33922;
squeal_samples[4239]=36008;
squeal_samples[4240]=38003;
squeal_samples[4241]=39912;
squeal_samples[4242]=41726;
squeal_samples[4243]=43473;
squeal_samples[4244]=45130;
squeal_samples[4245]=46719;
squeal_samples[4246]=48235;
squeal_samples[4247]=49684;
squeal_samples[4248]=51077;
squeal_samples[4249]=49887;
squeal_samples[4250]=44894;
squeal_samples[4251]=40160;
squeal_samples[4252]=35744;
squeal_samples[4253]=31601;
squeal_samples[4254]=27731;
squeal_samples[4255]=24110;
squeal_samples[4256]=20712;
squeal_samples[4257]=17545;
squeal_samples[4258]=14575;
squeal_samples[4259]=11807;
squeal_samples[4260]=9207;
squeal_samples[4261]=7880;
squeal_samples[4262]=10707;
squeal_samples[4263]=13801;
squeal_samples[4264]=16764;
squeal_samples[4265]=19607;
squeal_samples[4266]=22321;
squeal_samples[4267]=24920;
squeal_samples[4268]=27404;
squeal_samples[4269]=29771;
squeal_samples[4270]=32045;
squeal_samples[4271]=34214;
squeal_samples[4272]=36286;
squeal_samples[4273]=38271;
squeal_samples[4274]=40159;
squeal_samples[4275]=41973;
squeal_samples[4276]=43701;
squeal_samples[4277]=45353;
squeal_samples[4278]=46928;
squeal_samples[4279]=48438;
squeal_samples[4280]=49874;
squeal_samples[4281]=51252;
squeal_samples[4282]=49307;
squeal_samples[4283]=44296;
squeal_samples[4284]=39600;
squeal_samples[4285]=35219;
squeal_samples[4286]=31106;
squeal_samples[4287]=27273;
squeal_samples[4288]=23671;
squeal_samples[4289]=20310;
squeal_samples[4290]=17167;
squeal_samples[4291]=14220;
squeal_samples[4292]=11469;
squeal_samples[4293]=8893;
squeal_samples[4294]=8069;
squeal_samples[4295]=11097;
squeal_samples[4296]=14177;
squeal_samples[4297]=17123;
squeal_samples[4298]=19944;
squeal_samples[4299]=22652;
squeal_samples[4300]=25232;
squeal_samples[4301]=27705;
squeal_samples[4302]=30060;
squeal_samples[4303]=32315;
squeal_samples[4304]=34475;
squeal_samples[4305]=36533;
squeal_samples[4306]=38505;
squeal_samples[4307]=40390;
squeal_samples[4308]=42183;
squeal_samples[4309]=43902;
squeal_samples[4310]=45545;
squeal_samples[4311]=47112;
squeal_samples[4312]=48608;
squeal_samples[4313]=50048;
squeal_samples[4314]=51357;
squeal_samples[4315]=48652;
squeal_samples[4316]=43682;
squeal_samples[4317]=39026;
squeal_samples[4318]=34680;
squeal_samples[4319]=30604;
squeal_samples[4320]=26796;
squeal_samples[4321]=23232;
squeal_samples[4322]=19894;
squeal_samples[4323]=16773;
squeal_samples[4324]=13856;
squeal_samples[4325]=11127;
squeal_samples[4326]=8578;
squeal_samples[4327]=8332;
squeal_samples[4328]=11480;
squeal_samples[4329]=14540;
squeal_samples[4330]=17473;
squeal_samples[4331]=20280;
squeal_samples[4332]=22968;
squeal_samples[4333]=25536;
squeal_samples[4334]=27989;
squeal_samples[4335]=30334;
squeal_samples[4336]=32582;
squeal_samples[4337]=34724;
squeal_samples[4338]=36778;
squeal_samples[4339]=38730;
squeal_samples[4340]=40604;
squeal_samples[4341]=42394;
squeal_samples[4342]=44101;
squeal_samples[4343]=45731;
squeal_samples[4344]=47296;
squeal_samples[4345]=48780;
squeal_samples[4346]=50208;
squeal_samples[4347]=51362;
squeal_samples[4348]=47997;
squeal_samples[4349]=43070;
squeal_samples[4350]=38456;
squeal_samples[4351]=34138;
squeal_samples[4352]=30103;
squeal_samples[4353]=26327;
squeal_samples[4354]=22790;
squeal_samples[4355]=19478;
squeal_samples[4356]=16387;
squeal_samples[4357]=13494;
squeal_samples[4358]=10787;
squeal_samples[4359]=8257;
squeal_samples[4360]=8675;
squeal_samples[4361]=11861;
squeal_samples[4362]=14902;
squeal_samples[4363]=17815;
squeal_samples[4364]=20613;
squeal_samples[4365]=23276;
squeal_samples[4366]=25842;
squeal_samples[4367]=28277;
squeal_samples[4368]=30611;
squeal_samples[4369]=32838;
squeal_samples[4370]=34973;
squeal_samples[4371]=37013;
squeal_samples[4372]=38958;
squeal_samples[4373]=40816;
squeal_samples[4374]=42601;
squeal_samples[4375]=44297;
squeal_samples[4376]=45917;
squeal_samples[4377]=47470;
squeal_samples[4378]=48947;
squeal_samples[4379]=50370;
squeal_samples[4380]=51256;
squeal_samples[4381]=47355;
squeal_samples[4382]=42463;
squeal_samples[4383]=37888;
squeal_samples[4384]=33612;
squeal_samples[4385]=29597;
squeal_samples[4386]=25863;
squeal_samples[4387]=22348;
squeal_samples[4388]=19073;
squeal_samples[4389]=16001;
squeal_samples[4390]=13129;
squeal_samples[4391]=10449;
squeal_samples[4392]=7981;
squeal_samples[4393]=9072;
squeal_samples[4394]=12232;
squeal_samples[4395]=15258;
squeal_samples[4396]=18157;
squeal_samples[4397]=20940;
squeal_samples[4398]=23592;
squeal_samples[4399]=26135;
squeal_samples[4400]=28560;
squeal_samples[4401]=30878;
squeal_samples[4402]=33096;
squeal_samples[4403]=35224;
squeal_samples[4404]=37241;
squeal_samples[4405]=39186;
squeal_samples[4406]=41030;
squeal_samples[4407]=42804;
squeal_samples[4408]=44491;
squeal_samples[4409]=46105;
squeal_samples[4410]=47647;
squeal_samples[4411]=49120;
squeal_samples[4412]=50523;
squeal_samples[4413]=51051;
squeal_samples[4414]=46707;
squeal_samples[4415]=41868;
squeal_samples[4416]=37323;
squeal_samples[4417]=33083;
squeal_samples[4418]=29103;
squeal_samples[4419]=25397;
squeal_samples[4420]=21913;
squeal_samples[4421]=18662;
squeal_samples[4422]=15620;
squeal_samples[4423]=12773;
squeal_samples[4424]=10110;
squeal_samples[4425]=7799;
squeal_samples[4426]=9461;
squeal_samples[4427]=12605;
squeal_samples[4428]=15615;
squeal_samples[4429]=18501;
squeal_samples[4430]=21265;
squeal_samples[4431]=23903;
squeal_samples[4432]=26432;
squeal_samples[4433]=28844;
squeal_samples[4434]=31148;
squeal_samples[4435]=33357;
squeal_samples[4436]=35467;
squeal_samples[4437]=37481;
squeal_samples[4438]=39408;
squeal_samples[4439]=41247;
squeal_samples[4440]=43004;
squeal_samples[4441]=44683;
squeal_samples[4442]=46288;
squeal_samples[4443]=47817;
squeal_samples[4444]=49289;
squeal_samples[4445]=50681;
squeal_samples[4446]=50741;
squeal_samples[4447]=46070;
squeal_samples[4448]=41265;
squeal_samples[4449]=36765;
squeal_samples[4450]=32556;
squeal_samples[4451]=28620;
squeal_samples[4452]=24931;
squeal_samples[4453]=21484;
squeal_samples[4454]=18257;
squeal_samples[4455]=15236;
squeal_samples[4456]=12420;
squeal_samples[4457]=9775;
squeal_samples[4458]=7709;
squeal_samples[4459]=9847;
squeal_samples[4460]=12970;
squeal_samples[4461]=15972;
squeal_samples[4462]=18837;
squeal_samples[4463]=21586;
squeal_samples[4464]=24212;
squeal_samples[4465]=26727;
squeal_samples[4466]=29122;
squeal_samples[4467]=31414;
squeal_samples[4468]=33616;
squeal_samples[4469]=35709;
squeal_samples[4470]=37712;
squeal_samples[4471]=39629;
squeal_samples[4472]=41457;
squeal_samples[4473]=43206;
squeal_samples[4474]=44872;
squeal_samples[4475]=46470;
squeal_samples[4476]=47989;
squeal_samples[4477]=49449;
squeal_samples[4478]=50840;
squeal_samples[4479]=50328;
squeal_samples[4480]=45438;
squeal_samples[4481]=40676;
squeal_samples[4482]=36210;
squeal_samples[4483]=32032;
squeal_samples[4484]=28134;
squeal_samples[4485]=24478;
squeal_samples[4486]=21057;
squeal_samples[4487]=17854;
squeal_samples[4488]=14859;
squeal_samples[4489]=12064;
squeal_samples[4490]=9447;
squeal_samples[4491]=7701;
squeal_samples[4492]=10230;
squeal_samples[4493]=13344;
squeal_samples[4494]=16321;
squeal_samples[4495]=19179;
squeal_samples[4496]=21907;
squeal_samples[4497]=24522;
squeal_samples[4498]=27017;
squeal_samples[4499]=29400;
squeal_samples[4500]=31685;
squeal_samples[4501]=33869;
squeal_samples[4502]=35948;
squeal_samples[4503]=37948;
squeal_samples[4504]=39845;
squeal_samples[4505]=41669;
squeal_samples[4506]=43404;
squeal_samples[4507]=45064;
squeal_samples[4508]=46653;
squeal_samples[4509]=48167;
squeal_samples[4510]=49614;
squeal_samples[4511]=50997;
squeal_samples[4512]=49813;
squeal_samples[4513]=44813;
squeal_samples[4514]=40085;
squeal_samples[4515]=35660;
squeal_samples[4516]=31519;
squeal_samples[4517]=27649;
squeal_samples[4518]=24019;
squeal_samples[4519]=20632;
squeal_samples[4520]=17455;
squeal_samples[4521]=14487;
squeal_samples[4522]=11714;
squeal_samples[4523]=9117;
squeal_samples[4524]=7793;
squeal_samples[4525]=10614;
squeal_samples[4526]=13709;
squeal_samples[4527]=16675;
squeal_samples[4528]=19509;
squeal_samples[4529]=22229;
squeal_samples[4530]=24826;
squeal_samples[4531]=27309;
squeal_samples[4532]=29679;
squeal_samples[4533]=31951;
squeal_samples[4534]=34118;
squeal_samples[4535]=36194;
squeal_samples[4536]=38175;
squeal_samples[4537]=40067;
squeal_samples[4538]=41879;
squeal_samples[4539]=43599;
squeal_samples[4540]=45256;
squeal_samples[4541]=46827;
squeal_samples[4542]=48339;
squeal_samples[4543]=49775;
squeal_samples[4544]=51150;
squeal_samples[4545]=49965;
squeal_samples[4546]=44949;
squeal_samples[4547]=40216;
squeal_samples[4548]=35773;
squeal_samples[4549]=31629;
squeal_samples[4550]=27745;
squeal_samples[4551]=24118;
squeal_samples[4552]=20714;
squeal_samples[4553]=17541;
squeal_samples[4554]=14560;
squeal_samples[4555]=11781;
squeal_samples[4556]=9182;
squeal_samples[4557]=7847;
squeal_samples[4558]=10674;
squeal_samples[4559]=13760;
squeal_samples[4560]=16727;
squeal_samples[4561]=19555;
squeal_samples[4562]=22276;
squeal_samples[4563]=24866;
squeal_samples[4564]=27351;
squeal_samples[4565]=29715;
squeal_samples[4566]=31985;
squeal_samples[4567]=34149;
squeal_samples[4568]=36225;
squeal_samples[4569]=38204;
squeal_samples[4570]=40093;
squeal_samples[4571]=41902;
squeal_samples[4572]=43625;
squeal_samples[4573]=45275;
squeal_samples[4574]=46846;
squeal_samples[4575]=48359;
squeal_samples[4576]=49793;
squeal_samples[4577]=51170;
squeal_samples[4578]=49978;
squeal_samples[4579]=44965;
squeal_samples[4580]=40222;
squeal_samples[4581]=35790;
squeal_samples[4582]=31633;
squeal_samples[4583]=27759;
squeal_samples[4584]=24121;
squeal_samples[4585]=20723;
squeal_samples[4586]=17538;
squeal_samples[4587]=14568;
squeal_samples[4588]=11781;
squeal_samples[4589]=9187;
squeal_samples[4590]=7844;
squeal_samples[4591]=10671;
squeal_samples[4592]=13759;
squeal_samples[4593]=16723;
squeal_samples[4594]=19554;
squeal_samples[4595]=22273;
squeal_samples[4596]=24864;
squeal_samples[4597]=27349;
squeal_samples[4598]=29712;
squeal_samples[4599]=31976;
squeal_samples[4600]=34150;
squeal_samples[4601]=36214;
squeal_samples[4602]=38198;
squeal_samples[4603]=40084;
squeal_samples[4604]=41895;
squeal_samples[4605]=43618;
squeal_samples[4606]=45271;
squeal_samples[4607]=46845;
squeal_samples[4608]=48350;
squeal_samples[4609]=49786;
squeal_samples[4610]=51163;
squeal_samples[4611]=49968;
squeal_samples[4612]=44959;
squeal_samples[4613]=40213;
squeal_samples[4614]=35777;
squeal_samples[4615]=31627;
squeal_samples[4616]=27747;
squeal_samples[4617]=24114;
squeal_samples[4618]=20708;
squeal_samples[4619]=17531;
squeal_samples[4620]=14557;
squeal_samples[4621]=11774;
squeal_samples[4622]=9174;
squeal_samples[4623]=7836;
squeal_samples[4624]=10664;
squeal_samples[4625]=13744;
squeal_samples[4626]=16711;
squeal_samples[4627]=19541;
squeal_samples[4628]=22259;
squeal_samples[4629]=24852;
squeal_samples[4630]=27333;
squeal_samples[4631]=29702;
squeal_samples[4632]=31967;
squeal_samples[4633]=34136;
squeal_samples[4634]=36207;
squeal_samples[4635]=38184;
squeal_samples[4636]=40073;
squeal_samples[4637]=41879;
squeal_samples[4638]=43607;
squeal_samples[4639]=45256;
squeal_samples[4640]=46834;
squeal_samples[4641]=48334;
squeal_samples[4642]=49776;
squeal_samples[4643]=51147;
squeal_samples[4644]=49957;
squeal_samples[4645]=44946;
squeal_samples[4646]=40197;
squeal_samples[4647]=35774;
squeal_samples[4648]=31608;
squeal_samples[4649]=27741;
squeal_samples[4650]=24093;
squeal_samples[4651]=20702;
squeal_samples[4652]=17512;
squeal_samples[4653]=14547;
squeal_samples[4654]=11761;
squeal_samples[4655]=9158;
squeal_samples[4656]=7827;
squeal_samples[4657]=10645;
squeal_samples[4658]=13737;
squeal_samples[4659]=16693;
squeal_samples[4660]=19530;
squeal_samples[4661]=22245;
squeal_samples[4662]=24839;
squeal_samples[4663]=27321;
squeal_samples[4664]=29686;
squeal_samples[4665]=31957;
squeal_samples[4666]=34119;
squeal_samples[4667]=36198;
squeal_samples[4668]=38168;
squeal_samples[4669]=40065;
squeal_samples[4670]=41868;
squeal_samples[4671]=43591;
squeal_samples[4672]=45246;
squeal_samples[4673]=46818;
squeal_samples[4674]=48323;
squeal_samples[4675]=49761;
squeal_samples[4676]=51135;
squeal_samples[4677]=49944;
squeal_samples[4678]=44931;
squeal_samples[4679]=40188;
squeal_samples[4680]=35754;
squeal_samples[4681]=31602;
squeal_samples[4682]=27721;
squeal_samples[4683]=24085;
squeal_samples[4684]=20686;
squeal_samples[4685]=17500;
squeal_samples[4686]=14533;
squeal_samples[4687]=11747;
squeal_samples[4688]=9147;
squeal_samples[4689]=7812;
squeal_samples[4690]=10633;
squeal_samples[4691]=13724;
squeal_samples[4692]=16677;
squeal_samples[4693]=19523;
squeal_samples[4694]=22225;
squeal_samples[4695]=24831;
squeal_samples[4696]=27305;
squeal_samples[4697]=29674;
squeal_samples[4698]=31944;
squeal_samples[4699]=34107;
squeal_samples[4700]=36181;
squeal_samples[4701]=38159;
squeal_samples[4702]=40050;
squeal_samples[4703]=41855;
squeal_samples[4704]=43579;
squeal_samples[4705]=45231;
squeal_samples[4706]=46805;
squeal_samples[4707]=48312;
squeal_samples[4708]=49745;
squeal_samples[4709]=51124;
squeal_samples[4710]=49930;
squeal_samples[4711]=44917;
squeal_samples[4712]=40175;
squeal_samples[4713]=35743;
squeal_samples[4714]=31585;
squeal_samples[4715]=27713;
squeal_samples[4716]=24067;
squeal_samples[4717]=20675;
squeal_samples[4718]=17487;
squeal_samples[4719]=14518;
squeal_samples[4720]=11737;
squeal_samples[4721]=9130;
squeal_samples[4722]=7801;
squeal_samples[4723]=10621;
squeal_samples[4724]=13707;
squeal_samples[4725]=16669;
squeal_samples[4726]=19503;
squeal_samples[4727]=22219;
squeal_samples[4728]=24812;
squeal_samples[4729]=27296;
squeal_samples[4730]=29658;
squeal_samples[4731]=31931;
squeal_samples[4732]=34095;
squeal_samples[4733]=36167;
squeal_samples[4734]=38147;
squeal_samples[4735]=40034;
squeal_samples[4736]=41845;
squeal_samples[4737]=43561;
squeal_samples[4738]=45223;
squeal_samples[4739]=46790;
squeal_samples[4740]=48297;
squeal_samples[4741]=49735;
squeal_samples[4742]=51108;
squeal_samples[4743]=49917;
squeal_samples[4744]=44906;
squeal_samples[4745]=40160;
squeal_samples[4746]=35730;
squeal_samples[4747]=31573;
squeal_samples[4748]=27697;
squeal_samples[4749]=24057;
squeal_samples[4750]=20660;
squeal_samples[4751]=17475;
squeal_samples[4752]=14504;
squeal_samples[4753]=11725;
squeal_samples[4754]=9116;
squeal_samples[4755]=7788;
squeal_samples[4756]=10607;
squeal_samples[4757]=13696;
squeal_samples[4758]=16654;
squeal_samples[4759]=19492;
squeal_samples[4760]=22202;
squeal_samples[4761]=24804;
squeal_samples[4762]=27277;
squeal_samples[4763]=29651;
squeal_samples[4764]=31913;
squeal_samples[4765]=34084;
squeal_samples[4766]=36154;
squeal_samples[4767]=38132;
squeal_samples[4768]=40024;
squeal_samples[4769]=41828;
squeal_samples[4770]=43553;
squeal_samples[4771]=45204;
squeal_samples[4772]=46780;
squeal_samples[4773]=48284;
squeal_samples[4774]=49720;
squeal_samples[4775]=51096;
squeal_samples[4776]=49906;
squeal_samples[4777]=44888;
squeal_samples[4778]=40151;
squeal_samples[4779]=35714;
squeal_samples[4780]=31561;
squeal_samples[4781]=27684;
squeal_samples[4782]=24045;
squeal_samples[4783]=20643;
squeal_samples[4784]=17465;
squeal_samples[4785]=14490;
squeal_samples[4786]=11710;
squeal_samples[4787]=9106;
squeal_samples[4788]=7771;
squeal_samples[4789]=10597;
squeal_samples[4790]=13680;
squeal_samples[4791]=16644;
squeal_samples[4792]=19474;
squeal_samples[4793]=22194;
squeal_samples[4794]=24786;
squeal_samples[4795]=27268;
squeal_samples[4796]=29633;
squeal_samples[4797]=31905;
squeal_samples[4798]=34065;
squeal_samples[4799]=36147;
squeal_samples[4800]=38112;
squeal_samples[4801]=40017;
squeal_samples[4802]=41810;
squeal_samples[4803]=43543;
squeal_samples[4804]=45189;
squeal_samples[4805]=46767;
squeal_samples[4806]=48271;
squeal_samples[4807]=49707;
squeal_samples[4808]=51083;
squeal_samples[4809]=49892;
squeal_samples[4810]=44875;
squeal_samples[4811]=40139;
squeal_samples[4812]=35698;
squeal_samples[4813]=31552;
squeal_samples[4814]=27667;
squeal_samples[4815]=24033;
squeal_samples[4816]=20632;
squeal_samples[4817]=17448;
squeal_samples[4818]=14479;
squeal_samples[4819]=11696;
squeal_samples[4820]=9093;
squeal_samples[4821]=7759;
squeal_samples[4822]=10582;
squeal_samples[4823]=13667;
squeal_samples[4824]=16630;
squeal_samples[4825]=19463;
squeal_samples[4826]=22180;
squeal_samples[4827]=24772;
squeal_samples[4828]=27255;
squeal_samples[4829]=29621;
squeal_samples[4830]=31890;
squeal_samples[4831]=34055;
squeal_samples[4832]=36129;
squeal_samples[4833]=38104;
squeal_samples[4834]=40000;
squeal_samples[4835]=41799;
squeal_samples[4836]=43529;
squeal_samples[4837]=45176;
squeal_samples[4838]=46753;
squeal_samples[4839]=48260;
squeal_samples[4840]=49690;
squeal_samples[4841]=51074;
squeal_samples[4842]=49874;
squeal_samples[4843]=44866;
squeal_samples[4844]=40123;
squeal_samples[4845]=35686;
squeal_samples[4846]=31538;
squeal_samples[4847]=27653;
squeal_samples[4848]=24022;
squeal_samples[4849]=20616;
squeal_samples[4850]=17437;
squeal_samples[4851]=14465;
squeal_samples[4852]=11683;
squeal_samples[4853]=9079;
squeal_samples[4854]=7747;
squeal_samples[4855]=10567;
squeal_samples[4856]=13656;
squeal_samples[4857]=16616;
squeal_samples[4858]=19449;
squeal_samples[4859]=22166;
squeal_samples[4860]=24760;
squeal_samples[4861]=27241;
squeal_samples[4862]=29608;
squeal_samples[4863]=31877;
squeal_samples[4864]=34040;
squeal_samples[4865]=36118;
squeal_samples[4866]=38088;
squeal_samples[4867]=39988;
squeal_samples[4868]=41786;
squeal_samples[4869]=43514;
squeal_samples[4870]=45165;
squeal_samples[4871]=46737;
squeal_samples[4872]=48247;
squeal_samples[4873]=49677;
squeal_samples[4874]=51059;
squeal_samples[4875]=50520;
squeal_samples[4876]=45611;
squeal_samples[4877]=40827;
squeal_samples[4878]=36343;
squeal_samples[4879]=32152;
squeal_samples[4880]=28229;
squeal_samples[4881]=24553;
squeal_samples[4882]=21121;
squeal_samples[4883]=17907;
squeal_samples[4884]=14897;
squeal_samples[4885]=12087;
squeal_samples[4886]=9458;
squeal_samples[4887]=7705;
squeal_samples[4888]=10223;
squeal_samples[4889]=13334;
squeal_samples[4890]=16301;
squeal_samples[4891]=19157;
squeal_samples[4892]=21873;
squeal_samples[4893]=24488;
squeal_samples[4894]=26977;
squeal_samples[4895]=29356;
squeal_samples[4896]=31636;
squeal_samples[4897]=33811;
squeal_samples[4898]=35891;
squeal_samples[4899]=37876;
squeal_samples[4900]=39777;
squeal_samples[4901]=41595;
squeal_samples[4902]=43327;
squeal_samples[4903]=44983;
squeal_samples[4904]=46562;
squeal_samples[4905]=48082;
squeal_samples[4906]=49522;
squeal_samples[4907]=50905;
squeal_samples[4908]=50376;
squeal_samples[4909]=45480;
squeal_samples[4910]=40700;
squeal_samples[4911]=36219;
squeal_samples[4912]=32038;
squeal_samples[4913]=28116;
squeal_samples[4914]=24457;
squeal_samples[4915]=21017;
squeal_samples[4916]=17820;
squeal_samples[4917]=14811;
squeal_samples[4918]=12007;
squeal_samples[4919]=9382;
squeal_samples[4920]=7634;
squeal_samples[4921]=10155;
squeal_samples[4922]=13264;
squeal_samples[4923]=16244;
squeal_samples[4924]=19084;
squeal_samples[4925]=21821;
squeal_samples[4926]=24423;
squeal_samples[4927]=26922;
squeal_samples[4928]=29299;
squeal_samples[4929]=31578;
squeal_samples[4930]=33761;
squeal_samples[4931]=35839;
squeal_samples[4932]=37832;
squeal_samples[4933]=39729;
squeal_samples[4934]=41552;
squeal_samples[4935]=43277;
squeal_samples[4936]=44946;
squeal_samples[4937]=46520;
squeal_samples[4938]=48040;
squeal_samples[4939]=49483;
squeal_samples[4940]=50869;
squeal_samples[4941]=50899;
squeal_samples[4942]=46218;
squeal_samples[4943]=41385;
squeal_samples[4944]=36866;
squeal_samples[4945]=32636;
squeal_samples[4946]=28680;
squeal_samples[4947]=24978;
squeal_samples[4948]=21511;
squeal_samples[4949]=18274;
squeal_samples[4950]=15236;
squeal_samples[4951]=12408;
squeal_samples[4952]=9748;
squeal_samples[4953]=7676;
squeal_samples[4954]=9803;
squeal_samples[4955]=12927;
squeal_samples[4956]=15913;
squeal_samples[4957]=18779;
squeal_samples[4958]=21520;
squeal_samples[4959]=24136;
squeal_samples[4960]=26651;
squeal_samples[4961]=29034;
squeal_samples[4962]=31327;
squeal_samples[4963]=33520;
squeal_samples[4964]=35608;
squeal_samples[4965]=37611;
squeal_samples[4966]=39524;
squeal_samples[4967]=41343;
squeal_samples[4968]=43092;
squeal_samples[4969]=44752;
squeal_samples[4970]=46348;
squeal_samples[4971]=47867;
squeal_samples[4972]=49318;
squeal_samples[4973]=50708;
squeal_samples[4974]=51206;
squeal_samples[4975]=46854;
squeal_samples[4976]=41976;
squeal_samples[4977]=37421;
squeal_samples[4978]=33152;
squeal_samples[4979]=29163;
squeal_samples[4980]=25431;
squeal_samples[4981]=21934;
squeal_samples[4982]=18664;
squeal_samples[4983]=15607;
squeal_samples[4984]=12750;
squeal_samples[4985]=10074;
squeal_samples[4986]=7749;
squeal_samples[4987]=9398;
squeal_samples[4988]=12540;
squeal_samples[4989]=15544;
squeal_samples[4990]=18427;
squeal_samples[4991]=21177;
squeal_samples[4992]=23812;
squeal_samples[4993]=26337;
squeal_samples[4994]=28743;
squeal_samples[4995]=31045;
squeal_samples[4996]=33242;
squeal_samples[4997]=35350;
squeal_samples[4998]=37356;
squeal_samples[4999]=39283;
squeal_samples[5000]=41113;
squeal_samples[5001]=42871;
squeal_samples[5002]=44540;
squeal_samples[5003]=46144;
squeal_samples[5004]=47668;
squeal_samples[5005]=49133;
squeal_samples[5006]=50528;
squeal_samples[5007]=51404;
squeal_samples[5008]=47471;
squeal_samples[5009]=42561;
squeal_samples[5010]=37963;
squeal_samples[5011]=33662;
squeal_samples[5012]=29638;
squeal_samples[5013]=25874;
squeal_samples[5014]=22350;
squeal_samples[5015]=19053;
squeal_samples[5016]=15969;
squeal_samples[5017]=13082;
squeal_samples[5018]=10390;
squeal_samples[5019]=7908;
squeal_samples[5020]=8989;
squeal_samples[5021]=12145;
squeal_samples[5022]=15163;
squeal_samples[5023]=18059;
squeal_samples[5024]=20830;
squeal_samples[5025]=23475;
squeal_samples[5026]=26016;
squeal_samples[5027]=28432;
squeal_samples[5028]=30748;
squeal_samples[5029]=32960;
squeal_samples[5030]=35078;
squeal_samples[5031]=37102;
squeal_samples[5032]=39028;
squeal_samples[5033]=40881;
squeal_samples[5034]=42637;
squeal_samples[5035]=44328;
squeal_samples[5036]=45935;
squeal_samples[5037]=47469;
squeal_samples[5038]=48942;
squeal_samples[5039]=50343;
squeal_samples[5040]=51487;
squeal_samples[5041]=48090;
squeal_samples[5042]=43147;
squeal_samples[5043]=38509;
squeal_samples[5044]=34170;
squeal_samples[5045]=30114;
squeal_samples[5046]=26317;
squeal_samples[5047]=22764;
squeal_samples[5048]=19444;
squeal_samples[5049]=16329;
squeal_samples[5050]=13424;
squeal_samples[5051]=10702;
squeal_samples[5052]=8154;
squeal_samples[5053]=8576;
squeal_samples[5054]=11744;
squeal_samples[5055]=14782;
squeal_samples[5056]=17692;
squeal_samples[5057]=20473;
squeal_samples[5058]=23139;
squeal_samples[5059]=25691;
squeal_samples[5060]=28128;
squeal_samples[5061]=30450;
squeal_samples[5062]=32676;
squeal_samples[5063]=34805;
squeal_samples[5064]=36838;
squeal_samples[5065]=38784;
squeal_samples[5066]=40636;
squeal_samples[5067]=42416;
squeal_samples[5068]=44105;
squeal_samples[5069]=45728;
squeal_samples[5070]=47266;
squeal_samples[5071]=48749;
squeal_samples[5072]=50156;
squeal_samples[5073]=51466;
squeal_samples[5074]=48727;
squeal_samples[5075]=43735;
squeal_samples[5076]=39057;
squeal_samples[5077]=34682;
squeal_samples[5078]=30590;
squeal_samples[5079]=26766;
squeal_samples[5080]=23180;
squeal_samples[5081]=19832;
squeal_samples[5082]=16690;
squeal_samples[5083]=13759;
squeal_samples[5084]=11021;
squeal_samples[5085]=8451;
squeal_samples[5086]=8198;
squeal_samples[5087]=11339;
squeal_samples[5088]=14394;
squeal_samples[5089]=17321;
squeal_samples[5090]=20124;
squeal_samples[5091]=22799;
squeal_samples[5092]=25363;
squeal_samples[5093]=27816;
squeal_samples[5094]=30149;
squeal_samples[5095]=32393;
squeal_samples[5096]=34530;
squeal_samples[5097]=36576;
squeal_samples[5098]=38531;
squeal_samples[5099]=40396;
squeal_samples[5100]=42185;
squeal_samples[5101]=43881;
squeal_samples[5102]=45512;
squeal_samples[5103]=47071;
squeal_samples[5104]=48553;
squeal_samples[5105]=49973;
squeal_samples[5106]=51335;
squeal_samples[5107]=49361;
squeal_samples[5108]=44326;
squeal_samples[5109]=39612;
squeal_samples[5110]=35204;
squeal_samples[5111]=31075;
squeal_samples[5112]=27219;
squeal_samples[5113]=23603;
squeal_samples[5114]=20223;
squeal_samples[5115]=17061;
squeal_samples[5116]=14102;
squeal_samples[5117]=11339;
squeal_samples[5118]=8749;
squeal_samples[5119]=7912;
squeal_samples[5120]=10935;
squeal_samples[5121]=14006;
squeal_samples[5122]=16949;
squeal_samples[5123]=19763;
squeal_samples[5124]=22462;
squeal_samples[5125]=25033;
squeal_samples[5126]=27499;
squeal_samples[5127]=29850;
squeal_samples[5128]=32101;
squeal_samples[5129]=34257;
squeal_samples[5130]=36313;
squeal_samples[5131]=38279;
squeal_samples[5132]=40154;
squeal_samples[5133]=41951;
squeal_samples[5134]=43659;
squeal_samples[5135]=45301;
squeal_samples[5136]=46859;
squeal_samples[5137]=48362;
squeal_samples[5138]=49785;
squeal_samples[5139]=51153;
squeal_samples[5140]=49948;
squeal_samples[5141]=44924;
squeal_samples[5142]=40171;
squeal_samples[5143]=35728;
squeal_samples[5144]=31560;
squeal_samples[5145]=27676;
squeal_samples[5146]=24026;
squeal_samples[5147]=20622;
squeal_samples[5148]=17429;
squeal_samples[5149]=14450;
squeal_samples[5150]=11661;
squeal_samples[5151]=9052;
squeal_samples[5152]=7714;
squeal_samples[5153]=10531;
squeal_samples[5154]=13617;
squeal_samples[5155]=16573;
squeal_samples[5156]=19406;
squeal_samples[5157]=22118;
squeal_samples[5158]=24705;
squeal_samples[5159]=27189;
squeal_samples[5160]=29547;
squeal_samples[5161]=31817;
squeal_samples[5162]=33978;
squeal_samples[5163]=36044;
squeal_samples[5164]=38027;
squeal_samples[5165]=39910;
squeal_samples[5166]=41716;
squeal_samples[5167]=43439;
squeal_samples[5168]=45088;
squeal_samples[5169]=46658;
squeal_samples[5170]=48163;
squeal_samples[5171]=49600;
squeal_samples[5172]=50968;
squeal_samples[5173]=50442;
squeal_samples[5174]=45525;
squeal_samples[5175]=40733;
squeal_samples[5176]=36253;
squeal_samples[5177]=32053;
squeal_samples[5178]=28133;
squeal_samples[5179]=24461;
squeal_samples[5180]=21025;
squeal_samples[5181]=17801;
squeal_samples[5182]=14803;
squeal_samples[5183]=11983;
squeal_samples[5184]=9356;
squeal_samples[5185]=7602;
squeal_samples[5186]=10120;
squeal_samples[5187]=13225;
squeal_samples[5188]=16201;
squeal_samples[5189]=19046;
squeal_samples[5190]=21773;
squeal_samples[5191]=24377;
squeal_samples[5192]=26871;
squeal_samples[5193]=29247;
squeal_samples[5194]=31522;
squeal_samples[5195]=33698;
squeal_samples[5196]=35782;
squeal_samples[5197]=37769;
squeal_samples[5198]=39668;
squeal_samples[5199]=41482;
squeal_samples[5200]=43213;
squeal_samples[5201]=44869;
squeal_samples[5202]=46455;
squeal_samples[5203]=47965;
squeal_samples[5204]=49411;
squeal_samples[5205]=50788;
squeal_samples[5206]=50825;
squeal_samples[5207]=46135;
squeal_samples[5208]=41304;
squeal_samples[5209]=36780;
squeal_samples[5210]=32552;
squeal_samples[5211]=28597;
squeal_samples[5212]=24893;
squeal_samples[5213]=21424;
squeal_samples[5214]=18181;
squeal_samples[5215]=15150;
squeal_samples[5216]=12316;
squeal_samples[5217]=9660;
squeal_samples[5218]=7581;
squeal_samples[5219]=9708;
squeal_samples[5220]=12833;
squeal_samples[5221]=15816;
squeal_samples[5222]=18687;
squeal_samples[5223]=21422;
squeal_samples[5224]=24044;
squeal_samples[5225]=26555;
squeal_samples[5226]=28938;
squeal_samples[5227]=31234;
squeal_samples[5228]=33417;
squeal_samples[5229]=35514;
squeal_samples[5230]=37514;
squeal_samples[5231]=39417;
squeal_samples[5232]=41250;
squeal_samples[5233]=42984;
squeal_samples[5234]=44657;
squeal_samples[5235]=46246;
squeal_samples[5236]=47766;
squeal_samples[5237]=49218;
squeal_samples[5238]=50605;
squeal_samples[5239]=51473;
squeal_samples[5240]=47533;
squeal_samples[5241]=42612;
squeal_samples[5242]=38009;
squeal_samples[5243]=33690;
squeal_samples[5244]=29664;
squeal_samples[5245]=25886;
squeal_samples[5246]=22364;
squeal_samples[5247]=19051;
squeal_samples[5248]=15962;
squeal_samples[5249]=13075;
squeal_samples[5250]=10369;
squeal_samples[5251]=7893;
squeal_samples[5252]=8969;
squeal_samples[5253]=12113;
squeal_samples[5254]=15141;
squeal_samples[5255]=18023;
squeal_samples[5256]=20797;
squeal_samples[5257]=23440;
squeal_samples[5258]=25974;
squeal_samples[5259]=28396;
squeal_samples[5260]=30703;
squeal_samples[5261]=32917;
squeal_samples[5262]=35028;
squeal_samples[5263]=37049;
squeal_samples[5264]=38978;
squeal_samples[5265]=40825;
squeal_samples[5266]=42585;
squeal_samples[5267]=44266;
squeal_samples[5268]=45874;
squeal_samples[5269]=47412;
squeal_samples[5270]=48878;
squeal_samples[5271]=50281;
squeal_samples[5272]=51576;
squeal_samples[5273]=48824;
squeal_samples[5274]=43827;
squeal_samples[5275]=39138;
squeal_samples[5276]=34756;
squeal_samples[5277]=30652;
squeal_samples[5278]=26815;
squeal_samples[5279]=23228;
squeal_samples[5280]=19864;
squeal_samples[5281]=16722;
squeal_samples[5282]=13781;
squeal_samples[5283]=11033;
squeal_samples[5284]=8460;
squeal_samples[5285]=8200;
squeal_samples[5286]=11340;
squeal_samples[5287]=14394;
squeal_samples[5288]=17307;
squeal_samples[5289]=20115;
squeal_samples[5290]=22780;
squeal_samples[5291]=25354;
squeal_samples[5292]=27792;
squeal_samples[5293]=30132;
squeal_samples[5294]=32368;
squeal_samples[5295]=34503;
squeal_samples[5296]=36547;
squeal_samples[5297]=38499;
squeal_samples[5298]=40361;
squeal_samples[5299]=42149;
squeal_samples[5300]=43845;
squeal_samples[5301]=45476;
squeal_samples[5302]=47028;
squeal_samples[5303]=48512;
squeal_samples[5304]=49932;
squeal_samples[5305]=51287;
squeal_samples[5306]=50071;
squeal_samples[5307]=45033;
squeal_samples[5308]=40271;
squeal_samples[5309]=35816;
squeal_samples[5310]=31639;
squeal_samples[5311]=27746;
squeal_samples[5312]=24085;
squeal_samples[5313]=20674;
squeal_samples[5314]=17478;
squeal_samples[5315]=14486;
squeal_samples[5316]=11693;
squeal_samples[5317]=9079;
squeal_samples[5318]=7728;
squeal_samples[5319]=10546;
squeal_samples[5320]=13628;
squeal_samples[5321]=16582;
squeal_samples[5322]=19411;
squeal_samples[5323]=22118;
squeal_samples[5324]=24702;
squeal_samples[5325]=27183;
squeal_samples[5326]=29542;
squeal_samples[5327]=31804;
squeal_samples[5328]=33968;
squeal_samples[5329]=36030;
squeal_samples[5330]=38011;
squeal_samples[5331]=39891;
squeal_samples[5332]=41696;
squeal_samples[5333]=43414;
squeal_samples[5334]=45062;
squeal_samples[5335]=46633;
squeal_samples[5336]=48136;
squeal_samples[5337]=49570;
squeal_samples[5338]=50940;
squeal_samples[5339]=50969;
squeal_samples[5340]=46260;
squeal_samples[5341]=41426;
squeal_samples[5342]=36883;
squeal_samples[5343]=32647;
squeal_samples[5344]=28673;
squeal_samples[5345]=24972;
squeal_samples[5346]=21495;
squeal_samples[5347]=18242;
squeal_samples[5348]=15201;
squeal_samples[5349]=12359;
squeal_samples[5350]=9701;
squeal_samples[5351]=7615;
squeal_samples[5352]=9736;
squeal_samples[5353]=12861;
squeal_samples[5354]=15840;
squeal_samples[5355]=18703;
squeal_samples[5356]=21442;
squeal_samples[5357]=24056;
squeal_samples[5358]=26560;
squeal_samples[5359]=28948;
squeal_samples[5360]=31237;
squeal_samples[5361]=33428;
squeal_samples[5362]=35513;
squeal_samples[5363]=37511;
squeal_samples[5364]=39414;
squeal_samples[5365]=41244;
squeal_samples[5366]=42978;
squeal_samples[5367]=44645;
squeal_samples[5368]=46232;
squeal_samples[5369]=47751;
squeal_samples[5370]=49205;
squeal_samples[5371]=50589;
squeal_samples[5372]=51454;
squeal_samples[5373]=47510;
squeal_samples[5374]=42589;
squeal_samples[5375]=37982;
squeal_samples[5376]=33667;
squeal_samples[5377]=29637;
squeal_samples[5378]=25855;
squeal_samples[5379]=22332;
squeal_samples[5380]=19022;
squeal_samples[5381]=15930;
squeal_samples[5382]=13044;
squeal_samples[5383]=10335;
squeal_samples[5384]=7853;
squeal_samples[5385]=8931;
squeal_samples[5386]=12074;
squeal_samples[5387]=15101;
squeal_samples[5388]=17984;
squeal_samples[5389]=20759;
squeal_samples[5390]=23399;
squeal_samples[5391]=25936;
squeal_samples[5392]=28353;
squeal_samples[5393]=30660;
squeal_samples[5394]=32877;
squeal_samples[5395]=34986;
squeal_samples[5396]=37004;
squeal_samples[5397]=38942;
squeal_samples[5398]=40772;
squeal_samples[5399]=42548;
squeal_samples[5400]=44220;
squeal_samples[5401]=45836;
squeal_samples[5402]=47363;
squeal_samples[5403]=48831;
squeal_samples[5404]=50235;
squeal_samples[5405]=51525;
squeal_samples[5406]=48783;
squeal_samples[5407]=43774;
squeal_samples[5408]=39094;
squeal_samples[5409]=34704;
squeal_samples[5410]=30602;
squeal_samples[5411]=26772;
squeal_samples[5412]=23170;
squeal_samples[5413]=19817;
squeal_samples[5414]=16671;
squeal_samples[5415]=13731;
squeal_samples[5416]=10979;
squeal_samples[5417]=8414;
squeal_samples[5418]=8151;
squeal_samples[5419]=11291;
squeal_samples[5420]=14342;
squeal_samples[5421]=17265;
squeal_samples[5422]=20064;
squeal_samples[5423]=22736;
squeal_samples[5424]=25298;
squeal_samples[5425]=27743;
squeal_samples[5426]=30077;
squeal_samples[5427]=32316;
squeal_samples[5428]=34450;
squeal_samples[5429]=36502;
squeal_samples[5430]=38444;
squeal_samples[5431]=40317;
squeal_samples[5432]=42092;
squeal_samples[5433]=43796;
squeal_samples[5434]=45422;
squeal_samples[5435]=46977;
squeal_samples[5436]=48459;
squeal_samples[5437]=49878;
squeal_samples[5438]=51236;
squeal_samples[5439]=50018;
squeal_samples[5440]=44987;
squeal_samples[5441]=40218;
squeal_samples[5442]=35763;
squeal_samples[5443]=31587;
squeal_samples[5444]=27694;
squeal_samples[5445]=24038;
squeal_samples[5446]=20622;
squeal_samples[5447]=17424;
squeal_samples[5448]=14436;
squeal_samples[5449]=11638;
squeal_samples[5450]=9030;
squeal_samples[5451]=7673;
squeal_samples[5452]=10495;
squeal_samples[5453]=13575;
squeal_samples[5454]=16530;
squeal_samples[5455]=19359;
squeal_samples[5456]=22069;
squeal_samples[5457]=24652;
squeal_samples[5458]=27130;
squeal_samples[5459]=29489;
squeal_samples[5460]=31752;
squeal_samples[5461]=33913;
squeal_samples[5462]=35981;
squeal_samples[5463]=37958;
squeal_samples[5464]=39838;
squeal_samples[5465]=41643;
squeal_samples[5466]=43363;
squeal_samples[5467]=45006;
squeal_samples[5468]=46586;
squeal_samples[5469]=48080;
squeal_samples[5470]=49519;
squeal_samples[5471]=50889;
squeal_samples[5472]=50912;
squeal_samples[5473]=46214;
squeal_samples[5474]=41367;
squeal_samples[5475]=36837;
squeal_samples[5476]=32590;
squeal_samples[5477]=28629;
squeal_samples[5478]=24918;
squeal_samples[5479]=21443;
squeal_samples[5480]=18190;
squeal_samples[5481]=15148;
squeal_samples[5482]=12308;
squeal_samples[5483]=9648;
squeal_samples[5484]=7561;
squeal_samples[5485]=9687;
squeal_samples[5486]=12805;
squeal_samples[5487]=15797;
squeal_samples[5488]=18648;
squeal_samples[5489]=21391;
squeal_samples[5490]=24003;
squeal_samples[5491]=26508;
squeal_samples[5492]=28894;
squeal_samples[5493]=31189;
squeal_samples[5494]=33370;
squeal_samples[5495]=35466;
squeal_samples[5496]=37454;
squeal_samples[5497]=39365;
squeal_samples[5498]=41190;
squeal_samples[5499]=42925;
squeal_samples[5500]=44594;
squeal_samples[5501]=46184;
squeal_samples[5502]=47700;
squeal_samples[5503]=49152;
squeal_samples[5504]=50536;
squeal_samples[5505]=51403;
squeal_samples[5506]=47456;
squeal_samples[5507]=42539;
squeal_samples[5508]=37926;
squeal_samples[5509]=33619;
squeal_samples[5510]=29580;
squeal_samples[5511]=25807;
squeal_samples[5512]=22277;
squeal_samples[5513]=18970;
squeal_samples[5514]=15878;
squeal_samples[5515]=12991;
squeal_samples[5516]=10283;
squeal_samples[5517]=7802;
squeal_samples[5518]=8875;
squeal_samples[5519]=12027;
squeal_samples[5520]=15042;
squeal_samples[5521]=17939;
squeal_samples[5522]=20700;
squeal_samples[5523]=23352;
squeal_samples[5524]=25880;
squeal_samples[5525]=28303;
squeal_samples[5526]=30607;
squeal_samples[5527]=32825;
squeal_samples[5528]=34932;
squeal_samples[5529]=36955;
squeal_samples[5530]=38885;
squeal_samples[5531]=40726;
squeal_samples[5532]=42490;
squeal_samples[5533]=44172;
squeal_samples[5534]=45782;
squeal_samples[5535]=47308;
squeal_samples[5536]=48784;
squeal_samples[5537]=50178;
squeal_samples[5538]=51477;
squeal_samples[5539]=48727;
squeal_samples[5540]=43724;
squeal_samples[5541]=39041;
squeal_samples[5542]=34651;
squeal_samples[5543]=30551;
squeal_samples[5544]=26718;
squeal_samples[5545]=23120;
squeal_samples[5546]=19763;
squeal_samples[5547]=16619;
squeal_samples[5548]=13678;
squeal_samples[5549]=10928;
squeal_samples[5550]=8360;
squeal_samples[5551]=8101;
squeal_samples[5552]=11236;
squeal_samples[5553]=14291;
squeal_samples[5554]=17214;
squeal_samples[5555]=20008;
squeal_samples[5556]=22688;
squeal_samples[5557]=25242;
squeal_samples[5558]=27692;
squeal_samples[5559]=30026;
squeal_samples[5560]=32262;
squeal_samples[5561]=34399;
squeal_samples[5562]=36447;
squeal_samples[5563]=38395;
squeal_samples[5564]=40260;
squeal_samples[5565]=42046;
squeal_samples[5566]=43737;
squeal_samples[5567]=45374;
squeal_samples[5568]=46921;
squeal_samples[5569]=48409;
squeal_samples[5570]=49824;
squeal_samples[5571]=51183;
squeal_samples[5572]=50628;
squeal_samples[5573]=45695;
squeal_samples[5574]=40883;
squeal_samples[5575]=36384;
squeal_samples[5576]=32164;
squeal_samples[5577]=28228;
squeal_samples[5578]=24534;
squeal_samples[5579]=21084;
squeal_samples[5580]=17853;
squeal_samples[5581]=14830;
squeal_samples[5582]=12007;
squeal_samples[5583]=9366;
squeal_samples[5584]=7600;
squeal_samples[5585]=10118;
squeal_samples[5586]=13210;
squeal_samples[5587]=16180;
squeal_samples[5588]=19018;
squeal_samples[5589]=21741;
squeal_samples[5590]=24338;
squeal_samples[5591]=26827;
squeal_samples[5592]=29199;
squeal_samples[5593]=31471;
squeal_samples[5594]=33645;
squeal_samples[5595]=35720;
squeal_samples[5596]=37704;
squeal_samples[5597]=39599;
squeal_samples[5598]=41408;
squeal_samples[5599]=43139;
squeal_samples[5600]=44789;
squeal_samples[5601]=46370;
squeal_samples[5602]=47876;
squeal_samples[5603]=49319;
squeal_samples[5604]=50693;
squeal_samples[5605]=51546;
squeal_samples[5606]=47598;
squeal_samples[5607]=42661;
squeal_samples[5608]=38040;
squeal_samples[5609]=33724;
squeal_samples[5610]=29677;
squeal_samples[5611]=25898;
squeal_samples[5612]=22357;
squeal_samples[5613]=19046;
squeal_samples[5614]=15940;
squeal_samples[5615]=13050;
squeal_samples[5616]=10334;
squeal_samples[5617]=7846;
squeal_samples[5618]=8917;
squeal_samples[5619]=12063;
squeal_samples[5620]=15079;
squeal_samples[5621]=17969;
squeal_samples[5622]=20731;
squeal_samples[5623]=23381;
squeal_samples[5624]=25896;
squeal_samples[5625]=28327;
squeal_samples[5626]=30624;
squeal_samples[5627]=32841;
squeal_samples[5628]=34949;
squeal_samples[5629]=36961;
squeal_samples[5630]=38893;
squeal_samples[5631]=40731;
squeal_samples[5632]=42497;
squeal_samples[5633]=44169;
squeal_samples[5634]=45780;
squeal_samples[5635]=47309;
squeal_samples[5636]=48779;
squeal_samples[5637]=50178;
squeal_samples[5638]=51523;
squeal_samples[5639]=49525;
squeal_samples[5640]=44467;
squeal_samples[5641]=39728;
squeal_samples[5642]=35297;
squeal_samples[5643]=31152;
squeal_samples[5644]=27276;
squeal_samples[5645]=23646;
squeal_samples[5646]=20248;
squeal_samples[5647]=17071;
squeal_samples[5648]=14099;
squeal_samples[5649]=11317;
squeal_samples[5650]=8720;
squeal_samples[5651]=7868;
squeal_samples[5652]=10890;
squeal_samples[5653]=13950;
squeal_samples[5654]=16888;
squeal_samples[5655]=19696;
squeal_samples[5656]=22390;
squeal_samples[5657]=24951;
squeal_samples[5658]=27416;
squeal_samples[5659]=29756;
squeal_samples[5660]=32007;
squeal_samples[5661]=34154;
squeal_samples[5662]=36206;
squeal_samples[5663]=38165;
squeal_samples[5664]=40039;
squeal_samples[5665]=41828;
squeal_samples[5666]=43542;
squeal_samples[5667]=45170;
squeal_samples[5668]=46735;
squeal_samples[5669]=48220;
squeal_samples[5670]=49649;
squeal_samples[5671]=51014;
squeal_samples[5672]=51023;
squeal_samples[5673]=46313;
squeal_samples[5674]=41459;
squeal_samples[5675]=36913;
squeal_samples[5676]=32659;
squeal_samples[5677]=28687;
squeal_samples[5678]=24963;
squeal_samples[5679]=21485;
squeal_samples[5680]=18224;
squeal_samples[5681]=15179;
squeal_samples[5682]=12326;
squeal_samples[5683]=9663;
squeal_samples[5684]=7569;
squeal_samples[5685]=9689;
squeal_samples[5686]=12804;
squeal_samples[5687]=15787;
squeal_samples[5688]=18642;
squeal_samples[5689]=21381;
squeal_samples[5690]=23992;
squeal_samples[5691]=26492;
squeal_samples[5692]=28879;
squeal_samples[5693]=31159;
squeal_samples[5694]=33351;
squeal_samples[5695]=35434;
squeal_samples[5696]=37429;
squeal_samples[5697]=39337;
squeal_samples[5698]=41152;
squeal_samples[5699]=42899;
squeal_samples[5700]=44556;
squeal_samples[5701]=46144;
squeal_samples[5702]=47659;
squeal_samples[5703]=49110;
squeal_samples[5704]=50493;
squeal_samples[5705]=51607;
squeal_samples[5706]=48203;
squeal_samples[5707]=43227;
squeal_samples[5708]=38570;
squeal_samples[5709]=34208;
squeal_samples[5710]=30135;
squeal_samples[5711]=26319;
squeal_samples[5712]=22748;
squeal_samples[5713]=19405;
squeal_samples[5714]=16287;
squeal_samples[5715]=13358;
squeal_samples[5716]=10632;
squeal_samples[5717]=8071;
squeal_samples[5718]=8474;
squeal_samples[5719]=11640;
squeal_samples[5720]=14670;
squeal_samples[5721]=17577;
squeal_samples[5722]=20358;
squeal_samples[5723]=23010;
squeal_samples[5724]=25560;
squeal_samples[5725]=27989;
squeal_samples[5726]=30307;
squeal_samples[5727]=32529;
squeal_samples[5728]=34648;
squeal_samples[5729]=36680;
squeal_samples[5730]=38618;
squeal_samples[5731]=40466;
squeal_samples[5732]=42240;
squeal_samples[5733]=43923;
squeal_samples[5734]=45547;
squeal_samples[5735]=47084;
squeal_samples[5736]=48560;
squeal_samples[5737]=49967;
squeal_samples[5738]=51317;
squeal_samples[5739]=50094;
squeal_samples[5740]=45038;
squeal_samples[5741]=40268;
squeal_samples[5742]=35798;
squeal_samples[5743]=31620;
squeal_samples[5744]=27709;
squeal_samples[5745]=24047;
squeal_samples[5746]=20622;
squeal_samples[5747]=17417;
squeal_samples[5748]=14419;
squeal_samples[5749]=11620;
squeal_samples[5750]=9002;
squeal_samples[5751]=7644;
squeal_samples[5752]=10459;
squeal_samples[5753]=13538;
squeal_samples[5754]=16487;
squeal_samples[5755]=19314;
squeal_samples[5756]=22014;
squeal_samples[5757]=24603;
squeal_samples[5758]=27074;
squeal_samples[5759]=29432;
squeal_samples[5760]=31695;
squeal_samples[5761]=33855;
squeal_samples[5762]=35918;
squeal_samples[5763]=37887;
squeal_samples[5764]=39771;
squeal_samples[5765]=41574;
squeal_samples[5766]=43287;
squeal_samples[5767]=44936;
squeal_samples[5768]=46501;
squeal_samples[5769]=48004;
squeal_samples[5770]=49431;
squeal_samples[5771]=50805;
squeal_samples[5772]=51287;
squeal_samples[5773]=46907;
squeal_samples[5774]=42005;
squeal_samples[5775]=37428;
squeal_samples[5776]=33144;
squeal_samples[5777]=29127;
squeal_samples[5778]=25383;
squeal_samples[5779]=21868;
squeal_samples[5780]=18583;
squeal_samples[5781]=15508;
squeal_samples[5782]=12636;
squeal_samples[5783]=9948;
squeal_samples[5784]=7614;
squeal_samples[5785]=9251;
squeal_samples[5786]=12386;
squeal_samples[5787]=15384;
squeal_samples[5788]=18254;
squeal_samples[5789]=21009;
squeal_samples[5790]=23626;
squeal_samples[5791]=26151;
squeal_samples[5792]=28540;
squeal_samples[5793]=30849;
squeal_samples[5794]=33038;
squeal_samples[5795]=35140;
squeal_samples[5796]=37146;
squeal_samples[5797]=39065;
squeal_samples[5798]=40890;
squeal_samples[5799]=42644;
squeal_samples[5800]=44310;
squeal_samples[5801]=45910;
squeal_samples[5802]=47436;
squeal_samples[5803]=48889;
squeal_samples[5804]=50288;
squeal_samples[5805]=51561;
squeal_samples[5806]=48811;
squeal_samples[5807]=43793;
squeal_samples[5808]=39097;
squeal_samples[5809]=34701;
squeal_samples[5810]=30587;
squeal_samples[5811]=26743;
squeal_samples[5812]=23142;
squeal_samples[5813]=19776;
squeal_samples[5814]=16625;
squeal_samples[5815]=13676;
squeal_samples[5816]=10922;
squeal_samples[5817]=8342;
squeal_samples[5818]=8078;
squeal_samples[5819]=11214;
squeal_samples[5820]=14261;
squeal_samples[5821]=17182;
squeal_samples[5822]=19972;
squeal_samples[5823]=22652;
squeal_samples[5824]=25200;
squeal_samples[5825]=27655;
squeal_samples[5826]=29981;
squeal_samples[5827]=32214;
squeal_samples[5828]=34355;
squeal_samples[5829]=36386;
squeal_samples[5830]=38343;
squeal_samples[5831]=40199;
squeal_samples[5832]=41982;
squeal_samples[5833]=43681;
squeal_samples[5834]=45304;
squeal_samples[5835]=46857;
squeal_samples[5836]=48340;
squeal_samples[5837]=49755;
squeal_samples[5838]=51110;
squeal_samples[5839]=50557;
squeal_samples[5840]=45623;
squeal_samples[5841]=40806;
squeal_samples[5842]=36306;
squeal_samples[5843]=32084;
squeal_samples[5844]=28148;
squeal_samples[5845]=24454;
squeal_samples[5846]=21000;
squeal_samples[5847]=17770;
squeal_samples[5848]=14744;
squeal_samples[5849]=11918;
squeal_samples[5850]=9279;
squeal_samples[5851]=7507;
squeal_samples[5852]=10023;
squeal_samples[5853]=13118;
squeal_samples[5854]=16086;
squeal_samples[5855]=18926;
squeal_samples[5856]=21647;
squeal_samples[5857]=24246;
squeal_samples[5858]=26732;
squeal_samples[5859]=29105;
squeal_samples[5860]=31380;
squeal_samples[5861]=33550;
squeal_samples[5862]=35623;
squeal_samples[5863]=37611;
squeal_samples[5864]=39502;
squeal_samples[5865]=41314;
squeal_samples[5866]=43041;
squeal_samples[5867]=44696;
squeal_samples[5868]=46273;
squeal_samples[5869]=47779;
squeal_samples[5870]=49219;
squeal_samples[5871]=50595;
squeal_samples[5872]=51448;
squeal_samples[5873]=47500;
squeal_samples[5874]=42561;
squeal_samples[5875]=37941;
squeal_samples[5876]=33622;
squeal_samples[5877]=29571;
squeal_samples[5878]=25796;
squeal_samples[5879]=22251;
squeal_samples[5880]=18942;
squeal_samples[5881]=15843;
squeal_samples[5882]=12945;
squeal_samples[5883]=10230;
squeal_samples[5884]=7749;
squeal_samples[5885]=8815;
squeal_samples[5886]=11962;
squeal_samples[5887]=14973;
squeal_samples[5888]=17866;
squeal_samples[5889]=20629;
squeal_samples[5890]=23271;
squeal_samples[5891]=25805;
squeal_samples[5892]=28214;
squeal_samples[5893]=30529;
squeal_samples[5894]=32731;
squeal_samples[5895]=34846;
squeal_samples[5896]=36859;
squeal_samples[5897]=38789;
squeal_samples[5898]=40633;
squeal_samples[5899]=42388;
squeal_samples[5900]=44068;
squeal_samples[5901]=45674;
squeal_samples[5902]=47206;
squeal_samples[5903]=48672;
squeal_samples[5904]=50076;
squeal_samples[5905]=51416;
squeal_samples[5906]=50183;
squeal_samples[5907]=45124;
squeal_samples[5908]=40335;
squeal_samples[5909]=35859;
squeal_samples[5910]=31675;
squeal_samples[5911]=27755;
squeal_samples[5912]=24089;
squeal_samples[5913]=20651;
squeal_samples[5914]=17446;
squeal_samples[5915]=14440;
squeal_samples[5916]=11633;
squeal_samples[5917]=9005;
squeal_samples[5918]=7651;
squeal_samples[5919]=10458;
squeal_samples[5920]=13538;
squeal_samples[5921]=16485;
squeal_samples[5922]=19304;
squeal_samples[5923]=22013;
squeal_samples[5924]=24589;
squeal_samples[5925]=27059;
squeal_samples[5926]=29417;
squeal_samples[5927]=31671;
squeal_samples[5928]=33836;
squeal_samples[5929]=35893;
squeal_samples[5930]=37870;
squeal_samples[5931]=39740;
squeal_samples[5932]=41549;
squeal_samples[5933]=43260;
squeal_samples[5934]=44902;
squeal_samples[5935]=46471;
squeal_samples[5936]=47969;
squeal_samples[5937]=49401;
squeal_samples[5938]=50764;
squeal_samples[5939]=51254;
squeal_samples[5940]=46858;
squeal_samples[5941]=41966;
squeal_samples[5942]=37383;
squeal_samples[5943]=33095;
squeal_samples[5944]=29080;
squeal_samples[5945]=25333;
squeal_samples[5946]=21819;
squeal_samples[5947]=18536;
squeal_samples[5948]=15457;
squeal_samples[5949]=12589;
squeal_samples[5950]=9895;
squeal_samples[5951]=7556;
squeal_samples[5952]=9202;
squeal_samples[5953]=12328;
squeal_samples[5954]=15330;
squeal_samples[5955]=18204;
squeal_samples[5956]=20947;
squeal_samples[5957]=23581;
squeal_samples[5958]=26089;
squeal_samples[5959]=28491;
squeal_samples[5960]=30787;
squeal_samples[5961]=32984;
squeal_samples[5962]=35085;
squeal_samples[5963]=37088;
squeal_samples[5964]=39003;
squeal_samples[5965]=40833;
squeal_samples[5966]=42581;
squeal_samples[5967]=44253;
squeal_samples[5968]=45848;
squeal_samples[5969]=47378;
squeal_samples[5970]=48828;
squeal_samples[5971]=50228;
squeal_samples[5972]=51554;
squeal_samples[5973]=49558;
squeal_samples[5974]=44480;
squeal_samples[5975]=39741;
squeal_samples[5976]=35302;
squeal_samples[5977]=31140;
squeal_samples[5978]=27261;
squeal_samples[5979]=23618;
squeal_samples[5980]=20222;
squeal_samples[5981]=17034;
squeal_samples[5982]=14053;
squeal_samples[5983]=11278;
squeal_samples[5984]=8666;
squeal_samples[5985]=7813;
squeal_samples[5986]=10827;
squeal_samples[5987]=13889;
squeal_samples[5988]=16818;
squeal_samples[5989]=19632;
squeal_samples[5990]=22306;
squeal_samples[5991]=24888;
squeal_samples[5992]=27335;
squeal_samples[5993]=29683;
squeal_samples[5994]=31925;
squeal_samples[5995]=34072;
squeal_samples[5996]=36120;
squeal_samples[5997]=38079;
squeal_samples[5998]=39950;
squeal_samples[5999]=41738;
squeal_samples[6000]=43447;
squeal_samples[6001]=45075;
squeal_samples[6002]=46636;
squeal_samples[6003]=48122;
squeal_samples[6004]=49547;
squeal_samples[6005]=50907;
squeal_samples[6006]=51385;
squeal_samples[6007]=46984;
squeal_samples[6008]=42081;
squeal_samples[6009]=37487;
squeal_samples[6010]=33193;
squeal_samples[6011]=29174;
squeal_samples[6012]=25414;
squeal_samples[6013]=21894;
squeal_samples[6014]=18596;
squeal_samples[6015]=15525;
squeal_samples[6016]=12638;
squeal_samples[6017]=9947;
squeal_samples[6018]=7602;
squeal_samples[6019]=9243;
squeal_samples[6020]=12370;
squeal_samples[6021]=15368;
squeal_samples[6022]=18236;
squeal_samples[6023]=20979;
squeal_samples[6024]=23605;
squeal_samples[6025]=26121;
squeal_samples[6026]=28511;
squeal_samples[6027]=30811;
squeal_samples[6028]=33000;
squeal_samples[6029]=35104;
squeal_samples[6030]=37104;
squeal_samples[6031]=39017;
squeal_samples[6032]=40842;
squeal_samples[6033]=42595;
squeal_samples[6034]=44262;
squeal_samples[6035]=45859;
squeal_samples[6036]=47379;
squeal_samples[6037]=48841;
squeal_samples[6038]=50222;
squeal_samples[6039]=51561;
squeal_samples[6040]=49555;
squeal_samples[6041]=44482;
squeal_samples[6042]=39739;
squeal_samples[6043]=35293;
squeal_samples[6044]=31141;
squeal_samples[6045]=27252;
squeal_samples[6046]=23617;
squeal_samples[6047]=20212;
squeal_samples[6048]=17020;
squeal_samples[6049]=14049;
squeal_samples[6050]=11258;
squeal_samples[6051]=8656;
squeal_samples[6052]=7794;
squeal_samples[6053]=10813;
squeal_samples[6054]=13871;
squeal_samples[6055]=16809;
squeal_samples[6056]=19611;
squeal_samples[6057]=22296;
squeal_samples[6058]=24863;
squeal_samples[6059]=27321;
squeal_samples[6060]=29664;
squeal_samples[6061]=31908;
squeal_samples[6062]=34052;
squeal_samples[6063]=36106;
squeal_samples[6064]=38056;
squeal_samples[6065]=39932;
squeal_samples[6066]=41716;
squeal_samples[6067]=43426;
squeal_samples[6068]=45056;
squeal_samples[6069]=46614;
squeal_samples[6070]=48102;
squeal_samples[6071]=49527;
squeal_samples[6072]=50885;
squeal_samples[6073]=51365;
squeal_samples[6074]=46964;
squeal_samples[6075]=42059;
squeal_samples[6076]=37469;
squeal_samples[6077]=33170;
squeal_samples[6078]=29148;
squeal_samples[6079]=25390;
squeal_samples[6080]=21869;
squeal_samples[6081]=18582;
squeal_samples[6082]=15493;
squeal_samples[6083]=12616;
squeal_samples[6084]=9920;
squeal_samples[6085]=7579;
squeal_samples[6086]=9221;
squeal_samples[6087]=12345;
squeal_samples[6088]=15346;
squeal_samples[6089]=18207;
squeal_samples[6090]=20960;
squeal_samples[6091]=23578;
squeal_samples[6092]=26095;
squeal_samples[6093]=28491;
squeal_samples[6094]=30784;
squeal_samples[6095]=32982;
squeal_samples[6096]=35074;
squeal_samples[6097]=37083;
squeal_samples[6098]=38990;
squeal_samples[6099]=40829;
squeal_samples[6100]=42563;
squeal_samples[6101]=44240;
squeal_samples[6102]=45829;
squeal_samples[6103]=47356;
squeal_samples[6104]=48813;
squeal_samples[6105]=50204;
squeal_samples[6106]=51533;
squeal_samples[6107]=49529;
squeal_samples[6108]=44458;
squeal_samples[6109]=39709;
squeal_samples[6110]=35272;
squeal_samples[6111]=31111;
squeal_samples[6112]=27228;
squeal_samples[6113]=23591;
squeal_samples[6114]=20183;
squeal_samples[6115]=16999;
squeal_samples[6116]=14018;
squeal_samples[6117]=11236;
squeal_samples[6118]=8625;
squeal_samples[6119]=7777;
squeal_samples[6120]=10786;
squeal_samples[6121]=13846;
squeal_samples[6122]=16781;
squeal_samples[6123]=19585;
squeal_samples[6124]=22270;
squeal_samples[6125]=24838;
squeal_samples[6126]=27296;
squeal_samples[6127]=29636;
squeal_samples[6128]=31881;
squeal_samples[6129]=34029;
squeal_samples[6130]=36076;
squeal_samples[6131]=38035;
squeal_samples[6132]=39902;
squeal_samples[6133]=41692;
squeal_samples[6134]=43399;
squeal_samples[6135]=45031;
squeal_samples[6136]=46587;
squeal_samples[6137]=48076;
squeal_samples[6138]=49502;
squeal_samples[6139]=50858;
squeal_samples[6140]=51340;
squeal_samples[6141]=46937;
squeal_samples[6142]=42034;
squeal_samples[6143]=37441;
squeal_samples[6144]=33146;
squeal_samples[6145]=29121;
squeal_samples[6146]=25364;
squeal_samples[6147]=21844;
squeal_samples[6148]=18554;
squeal_samples[6149]=15468;
squeal_samples[6150]=12590;
squeal_samples[6151]=9893;
squeal_samples[6152]=7556;
squeal_samples[6153]=9190;
squeal_samples[6154]=12323;
squeal_samples[6155]=15318;
squeal_samples[6156]=18182;
squeal_samples[6157]=20933;
squeal_samples[6158]=23553;
squeal_samples[6159]=26067;
squeal_samples[6160]=28468;
squeal_samples[6161]=30755;
squeal_samples[6162]=32957;
squeal_samples[6163]=35049;
squeal_samples[6164]=37054;
squeal_samples[6165]=38968;
squeal_samples[6166]=40799;
squeal_samples[6167]=42539;
squeal_samples[6168]=44215;
squeal_samples[6169]=45801;
squeal_samples[6170]=47331;
squeal_samples[6171]=48786;
squeal_samples[6172]=50178;
squeal_samples[6173]=51508;
squeal_samples[6174]=49502;
squeal_samples[6175]=44433;
squeal_samples[6176]=39681;
squeal_samples[6177]=35248;
squeal_samples[6178]=31083;
squeal_samples[6179]=27203;
squeal_samples[6180]=23566;
squeal_samples[6181]=20155;
squeal_samples[6182]=16975;
squeal_samples[6183]=13991;
squeal_samples[6184]=11209;
squeal_samples[6185]=8602;
squeal_samples[6186]=7748;
squeal_samples[6187]=10762;
squeal_samples[6188]=13818;
squeal_samples[6189]=16757;
squeal_samples[6190]=19558;
squeal_samples[6191]=22245;
squeal_samples[6192]=24811;
squeal_samples[6193]=27269;
squeal_samples[6194]=29611;
squeal_samples[6195]=31856;
squeal_samples[6196]=34002;
squeal_samples[6197]=36050;
squeal_samples[6198]=38009;
squeal_samples[6199]=39875;
squeal_samples[6200]=41667;
squeal_samples[6201]=43373;
squeal_samples[6202]=45004;
squeal_samples[6203]=46561;
squeal_samples[6204]=48051;
squeal_samples[6205]=49474;
squeal_samples[6206]=50835;
squeal_samples[6207]=51310;
squeal_samples[6208]=46914;
squeal_samples[6209]=42006;
squeal_samples[6210]=37416;
squeal_samples[6211]=33121;
squeal_samples[6212]=29092;
squeal_samples[6213]=25341;
squeal_samples[6214]=21815;
squeal_samples[6215]=18531;
squeal_samples[6216]=15440;
squeal_samples[6217]=12564;
squeal_samples[6218]=9868;
squeal_samples[6219]=7528;
squeal_samples[6220]=9166;
squeal_samples[6221]=12297;
squeal_samples[6222]=15290;
squeal_samples[6223]=18157;
squeal_samples[6224]=20907;
squeal_samples[6225]=23526;
squeal_samples[6226]=26042;
squeal_samples[6227]=28441;
squeal_samples[6228]=30730;
squeal_samples[6229]=32930;
squeal_samples[6230]=35024;
squeal_samples[6231]=37025;
squeal_samples[6232]=38945;
squeal_samples[6233]=40770;
squeal_samples[6234]=42515;
squeal_samples[6235]=44187;
squeal_samples[6236]=45775;
squeal_samples[6237]=47307;
squeal_samples[6238]=48755;
squeal_samples[6239]=50155;
squeal_samples[6240]=51479;
squeal_samples[6241]=50238;
squeal_samples[6242]=45166;
squeal_samples[6243]=40369;
squeal_samples[6244]=35881;
squeal_samples[6245]=31684;
squeal_samples[6246]=27757;
squeal_samples[6247]=24081;
squeal_samples[6248]=20642;
squeal_samples[6249]=17425;
squeal_samples[6250]=14410;
squeal_samples[6251]=11602;
squeal_samples[6252]=8966;
squeal_samples[6253]=7603;
squeal_samples[6254]=10408;
squeal_samples[6255]=13484;
squeal_samples[6256]=16429;
squeal_samples[6257]=19247;
squeal_samples[6258]=21946;
squeal_samples[6259]=24524;
squeal_samples[6260]=26993;
squeal_samples[6261]=29346;
squeal_samples[6262]=31602;
squeal_samples[6263]=33759;
squeal_samples[6264]=35812;
squeal_samples[6265]=37786;
squeal_samples[6266]=39661;
squeal_samples[6267]=41460;
squeal_samples[6268]=43174;
squeal_samples[6269]=44814;
squeal_samples[6270]=46378;
squeal_samples[6271]=47878;
squeal_samples[6272]=49306;
squeal_samples[6273]=50673;
squeal_samples[6274]=51513;
squeal_samples[6275]=47549;
squeal_samples[6276]=42600;
squeal_samples[6277]=37965;
squeal_samples[6278]=33632;
squeal_samples[6279]=29579;
squeal_samples[6280]=25790;
squeal_samples[6281]=22236;
squeal_samples[6282]=18916;
squeal_samples[6283]=15805;
squeal_samples[6284]=12903;
squeal_samples[6285]=10182;
squeal_samples[6286]=7690;
squeal_samples[6287]=8751;
squeal_samples[6288]=11898;
squeal_samples[6289]=14903;
squeal_samples[6290]=17791;
squeal_samples[6291]=20553;
squeal_samples[6292]=23192;
squeal_samples[6293]=25717;
squeal_samples[6294]=28132;
squeal_samples[6295]=30432;
squeal_samples[6296]=32645;
squeal_samples[6297]=34745;
squeal_samples[6298]=36765;
squeal_samples[6299]=38685;
squeal_samples[6300]=40533;
squeal_samples[6301]=42277;
squeal_samples[6302]=43963;
squeal_samples[6303]=45563;
squeal_samples[6304]=47101;
squeal_samples[6305]=48557;
squeal_samples[6306]=49960;
squeal_samples[6307]=51291;
squeal_samples[6308]=50728;
squeal_samples[6309]=45761;
squeal_samples[6310]=40931;
squeal_samples[6311]=36403;
squeal_samples[6312]=32168;
squeal_samples[6313]=28214;
squeal_samples[6314]=24506;
squeal_samples[6315]=21034;
squeal_samples[6316]=17788;
squeal_samples[6317]=14756;
squeal_samples[6318]=11916;
squeal_samples[6319]=9262;
squeal_samples[6320]=7483;
squeal_samples[6321]=9992;
squeal_samples[6322]=13082;
squeal_samples[6323]=16045;
squeal_samples[6324]=18878;
squeal_samples[6325]=21588;
squeal_samples[6326]=24184;
squeal_samples[6327]=26664;
squeal_samples[6328]=29030;
squeal_samples[6329]=31300;
squeal_samples[6330]=33464;
squeal_samples[6331]=35540;
squeal_samples[6332]=37513;
squeal_samples[6333]=39409;
squeal_samples[6334]=41214;
squeal_samples[6335]=42938;
squeal_samples[6336]=44585;
squeal_samples[6337]=46163;
squeal_samples[6338]=47666;
squeal_samples[6339]=49100;
squeal_samples[6340]=50478;
squeal_samples[6341]=51739;
squeal_samples[6342]=48966;
squeal_samples[6343]=43919;
squeal_samples[6344]=39206;
squeal_samples[6345]=34787;
squeal_samples[6346]=30657;
squeal_samples[6347]=26794;
squeal_samples[6348]=23179;
squeal_samples[6349]=19792;
squeal_samples[6350]=16630;
squeal_samples[6351]=13667;
squeal_samples[6352]=10898;
squeal_samples[6353]=8307;
squeal_samples[6354]=8031;
squeal_samples[6355]=11163;
squeal_samples[6356]=14206;
squeal_samples[6357]=17116;
squeal_samples[6358]=19903;
squeal_samples[6359]=22574;
squeal_samples[6360]=25126;
squeal_samples[6361]=27563;
squeal_samples[6362]=29891;
squeal_samples[6363]=32117;
squeal_samples[6364]=34250;
squeal_samples[6365]=36284;
squeal_samples[6366]=38230;
squeal_samples[6367]=40082;
squeal_samples[6368]=41861;
squeal_samples[6369]=43557;
squeal_samples[6370]=45177;
squeal_samples[6371]=46724;
squeal_samples[6372]=48202;
squeal_samples[6373]=49614;
squeal_samples[6374]=50972;
squeal_samples[6375]=51432;
squeal_samples[6376]=47025;
squeal_samples[6377]=42099;
squeal_samples[6378]=37506;
squeal_samples[6379]=33193;
squeal_samples[6380]=29167;
squeal_samples[6381]=25401;
squeal_samples[6382]=21872;
squeal_samples[6383]=18570;
squeal_samples[6384]=15487;
squeal_samples[6385]=12594;
squeal_samples[6386]=9896;
squeal_samples[6387]=7548;
squeal_samples[6388]=9181;
squeal_samples[6389]=12309;
squeal_samples[6390]=15299;
squeal_samples[6391]=18165;
squeal_samples[6392]=20903;
squeal_samples[6393]=23528;
squeal_samples[6394]=26040;
squeal_samples[6395]=28436;
squeal_samples[6396]=30724;
squeal_samples[6397]=32919;
squeal_samples[6398]=35011;
squeal_samples[6399]=37012;
squeal_samples[6400]=38919;
squeal_samples[6401]=40750;
squeal_samples[6402]=42493;
squeal_samples[6403]=44158;
squeal_samples[6404]=45755;
squeal_samples[6405]=47277;
squeal_samples[6406]=48724;
squeal_samples[6407]=50122;
squeal_samples[6408]=51445;
squeal_samples[6409]=50206;
squeal_samples[6410]=45127;
squeal_samples[6411]=40330;
squeal_samples[6412]=35843;
squeal_samples[6413]=31640;
squeal_samples[6414]=27713;
squeal_samples[6415]=24038;
squeal_samples[6416]=20592;
squeal_samples[6417]=17374;
squeal_samples[6418]=14364;
squeal_samples[6419]=11549;
squeal_samples[6420]=8916;
squeal_samples[6421]=7549;
squeal_samples[6422]=10363;
squeal_samples[6423]=13427;
squeal_samples[6424]=16375;
squeal_samples[6425]=19192;
squeal_samples[6426]=21890;
squeal_samples[6427]=24471;
squeal_samples[6428]=26938;
squeal_samples[6429]=29292;
squeal_samples[6430]=31546;
squeal_samples[6431]=33697;
squeal_samples[6432]=35761;
squeal_samples[6433]=37722;
squeal_samples[6434]=39605;
squeal_samples[6435]=41397;
squeal_samples[6436]=43114;
squeal_samples[6437]=44755;
squeal_samples[6438]=46317;
squeal_samples[6439]=47817;
squeal_samples[6440]=49247;
squeal_samples[6441]=50610;
squeal_samples[6442]=51709;
squeal_samples[6443]=48277;
squeal_samples[6444]=43279;
squeal_samples[6445]=38598;
squeal_samples[6446]=34225;
squeal_samples[6447]=30121;
squeal_samples[6448]=26294;
squeal_samples[6449]=22704;
squeal_samples[6450]=19348;
squeal_samples[6451]=16207;
squeal_samples[6452]=13279;
squeal_samples[6453]=10522;
squeal_samples[6454]=7962;
squeal_samples[6455]=8354;
squeal_samples[6456]=11515;
squeal_samples[6457]=14535;
squeal_samples[6458]=17438;
squeal_samples[6459]=20203;
squeal_samples[6460]=22863;
squeal_samples[6461]=25394;
squeal_samples[6462]=27822;
squeal_samples[6463]=30136;
squeal_samples[6464]=32353;
squeal_samples[6465]=34471;
squeal_samples[6466]=36496;
squeal_samples[6467]=38426;
squeal_samples[6468]=40276;
squeal_samples[6469]=42033;
squeal_samples[6470]=43729;
squeal_samples[6471]=45335;
squeal_samples[6472]=46876;
squeal_samples[6473]=48348;
squeal_samples[6474]=49747;
squeal_samples[6475]=51098;
squeal_samples[6476]=51087;
squeal_samples[6477]=46357;
squeal_samples[6478]=41472;
squeal_samples[6479]=36912;
squeal_samples[6480]=32640;
squeal_samples[6481]=28640;
squeal_samples[6482]=24911;
squeal_samples[6483]=21405;
squeal_samples[6484]=18137;
squeal_samples[6485]=15070;
squeal_samples[6486]=12210;
squeal_samples[6487]=9532;
squeal_samples[6488]=7426;
squeal_samples[6489]=9537;
squeal_samples[6490]=12649;
squeal_samples[6491]=15625;
squeal_samples[6492]=18476;
squeal_samples[6493]=21203;
squeal_samples[6494]=23808;
squeal_samples[6495]=26305;
squeal_samples[6496]=28684;
squeal_samples[6497]=30961;
squeal_samples[6498]=33146;
squeal_samples[6499]=35227;
squeal_samples[6500]=37216;
squeal_samples[6501]=39113;
squeal_samples[6502]=40935;
squeal_samples[6503]=42668;
squeal_samples[6504]=44328;
squeal_samples[6505]=45908;
squeal_samples[6506]=47425;
squeal_samples[6507]=48862;
squeal_samples[6508]=50252;
squeal_samples[6509]=51569;
squeal_samples[6510]=49558;
squeal_samples[6511]=44474;
squeal_samples[6512]=39715;
squeal_samples[6513]=35259;
squeal_samples[6514]=31098;
squeal_samples[6515]=27199;
squeal_samples[6516]=23555;
squeal_samples[6517]=20139;
squeal_samples[6518]=16950;
squeal_samples[6519]=13960;
squeal_samples[6520]=11168;
squeal_samples[6521]=8559;
squeal_samples[6522]=7698;
squeal_samples[6523]=10711;
squeal_samples[6524]=13766;
squeal_samples[6525]=16692;
squeal_samples[6526]=19502;
squeal_samples[6527]=22181;
squeal_samples[6528]=24747;
squeal_samples[6529]=27197;
squeal_samples[6530]=29539;
squeal_samples[6531]=31780;
squeal_samples[6532]=33924;
squeal_samples[6533]=35969;
squeal_samples[6534]=37925;
squeal_samples[6535]=39795;
squeal_samples[6536]=41582;
squeal_samples[6537]=43288;
squeal_samples[6538]=44912;
squeal_samples[6539]=46473;
squeal_samples[6540]=47953;
squeal_samples[6541]=49384;
squeal_samples[6542]=50732;
squeal_samples[6543]=51575;
squeal_samples[6544]=47593;
squeal_samples[6545]=42644;
squeal_samples[6546]=37995;
squeal_samples[6547]=33654;
squeal_samples[6548]=29593;
squeal_samples[6549]=25789;
squeal_samples[6550]=22238;
squeal_samples[6551]=18905;
squeal_samples[6552]=15795;
squeal_samples[6553]=12883;
squeal_samples[6554]=10160;
squeal_samples[6555]=7659;
squeal_samples[6556]=8718;
squeal_samples[6557]=11856;
squeal_samples[6558]=14866;
squeal_samples[6559]=17749;
squeal_samples[6560]=20503;
squeal_samples[6561]=23141;
squeal_samples[6562]=25667;
squeal_samples[6563]=28073;
squeal_samples[6564]=30381;
squeal_samples[6565]=32577;
squeal_samples[6566]=34690;
squeal_samples[6567]=36698;
squeal_samples[6568]=38623;
squeal_samples[6569]=40459;
squeal_samples[6570]=42218;
squeal_samples[6571]=43890;
squeal_samples[6572]=45494;
squeal_samples[6573]=47028;
squeal_samples[6574]=48482;
squeal_samples[6575]=49890;
squeal_samples[6576]=51213;
squeal_samples[6577]=50649;
squeal_samples[6578]=45683;
squeal_samples[6579]=40854;
squeal_samples[6580]=36319;
squeal_samples[6581]=32086;
squeal_samples[6582]=28124;
squeal_samples[6583]=24417;
squeal_samples[6584]=20946;
squeal_samples[6585]=17699;
squeal_samples[6586]=14663;
squeal_samples[6587]=11825;
squeal_samples[6588]=9170;
squeal_samples[6589]=7387;
squeal_samples[6590]=9899;
squeal_samples[6591]=12988;
squeal_samples[6592]=15950;
squeal_samples[6593]=18784;
squeal_samples[6594]=21494;
squeal_samples[6595]=24089;
squeal_samples[6596]=26570;
squeal_samples[6597]=28937;
squeal_samples[6598]=31204;
squeal_samples[6599]=33372;
squeal_samples[6600]=35438;
squeal_samples[6601]=37419;
squeal_samples[6602]=39310;
squeal_samples[6603]=41114;
squeal_samples[6604]=42843;
squeal_samples[6605]=44487;
squeal_samples[6606]=46061;
squeal_samples[6607]=47566;
squeal_samples[6608]=49001;
squeal_samples[6609]=50376;
squeal_samples[6610]=51690;
squeal_samples[6611]=49668;
squeal_samples[6612]=44577;
squeal_samples[6613]=39809;
squeal_samples[6614]=35347;
squeal_samples[6615]=31175;
squeal_samples[6616]=27270;
squeal_samples[6617]=23616;
squeal_samples[6618]=20200;
squeal_samples[6619]=17000;
squeal_samples[6620]=14009;
squeal_samples[6621]=11209;
squeal_samples[6622]=8594;
squeal_samples[6623]=7726;
squeal_samples[6624]=10734;
squeal_samples[6625]=13794;
squeal_samples[6626]=16714;
squeal_samples[6627]=19520;
squeal_samples[6628]=22192;
squeal_samples[6629]=24765;
squeal_samples[6630]=27203;
squeal_samples[6631]=29551;
squeal_samples[6632]=31787;
squeal_samples[6633]=33929;
squeal_samples[6634]=35972;
squeal_samples[6635]=37928;
squeal_samples[6636]=39794;
squeal_samples[6637]=41575;
squeal_samples[6638]=43279;
squeal_samples[6639]=44909;
squeal_samples[6640]=46459;
squeal_samples[6641]=47952;
squeal_samples[6642]=49366;
squeal_samples[6643]=50728;
squeal_samples[6644]=51814;
squeal_samples[6645]=48371;
squeal_samples[6646]=43363;
squeal_samples[6647]=38672;
squeal_samples[6648]=34285;
squeal_samples[6649]=30179;
squeal_samples[6650]=26339;
squeal_samples[6651]=22743;
squeal_samples[6652]=19385;
squeal_samples[6653]=16230;
squeal_samples[6654]=13291;
squeal_samples[6655]=10537;
squeal_samples[6656]=7968;
squeal_samples[6657]=8351;
squeal_samples[6658]=11513;
squeal_samples[6659]=14531;
squeal_samples[6660]=17423;
squeal_samples[6661]=20191;
squeal_samples[6662]=22846;
squeal_samples[6663]=25377;
squeal_samples[6664]=27802;
squeal_samples[6665]=30111;
squeal_samples[6666]=32321;
squeal_samples[6667]=34444;
squeal_samples[6668]=36461;
squeal_samples[6669]=38395;
squeal_samples[6670]=40235;
squeal_samples[6671]=42002;
squeal_samples[6672]=43689;
squeal_samples[6673]=45297;
squeal_samples[6674]=46832;
squeal_samples[6675]=48303;
squeal_samples[6676]=49699;
squeal_samples[6677]=51050;
squeal_samples[6678]=51499;
squeal_samples[6679]=47083;
squeal_samples[6680]=42153;
squeal_samples[6681]=37541;
squeal_samples[6682]=33223;
squeal_samples[6683]=29182;
squeal_samples[6684]=25409;
squeal_samples[6685]=21872;
squeal_samples[6686]=18562;
squeal_samples[6687]=15468;
squeal_samples[6688]=12576;
squeal_samples[6689]=9867;
squeal_samples[6690]=7512;
squeal_samples[6691]=9146;
squeal_samples[6692]=12262;
squeal_samples[6693]=15255;
squeal_samples[6694]=18113;
squeal_samples[6695]=20857;
squeal_samples[6696]=23474;
squeal_samples[6697]=25983;
squeal_samples[6698]=28368;
squeal_samples[6699]=30663;
squeal_samples[6700]=32852;
squeal_samples[6701]=34943;
squeal_samples[6702]=36941;
squeal_samples[6703]=38850;
squeal_samples[6704]=40674;
squeal_samples[6705]=42419;
squeal_samples[6706]=44081;
squeal_samples[6707]=45675;
squeal_samples[6708]=47195;
squeal_samples[6709]=48645;
squeal_samples[6710]=50034;
squeal_samples[6711]=51358;
squeal_samples[6712]=50779;
squeal_samples[6713]=45804;
squeal_samples[6714]=40958;
squeal_samples[6715]=36418;
squeal_samples[6716]=32179;
squeal_samples[6717]=28203;
squeal_samples[6718]=24488;
squeal_samples[6719]=21012;
squeal_samples[6720]=17760;
squeal_samples[6721]=14712;
squeal_samples[6722]=11866;
squeal_samples[6723]=9208;
squeal_samples[6724]=7423;
squeal_samples[6725]=9924;
squeal_samples[6726]=13014;
squeal_samples[6727]=15965;
squeal_samples[6728]=18804;
squeal_samples[6729]=21510;
squeal_samples[6730]=24102;
squeal_samples[6731]=26576;
squeal_samples[6732]=28944;
squeal_samples[6733]=31205;
squeal_samples[6734]=33374;
squeal_samples[6735]=35438;
squeal_samples[6736]=37419;
squeal_samples[6737]=39299;
squeal_samples[6738]=41111;
squeal_samples[6739]=42823;
squeal_samples[6740]=44481;
squeal_samples[6741]=46045;
squeal_samples[6742]=47551;
squeal_samples[6743]=48986;
squeal_samples[6744]=50356;
squeal_samples[6745]=51670;
squeal_samples[6746]=49642;
squeal_samples[6747]=44551;
squeal_samples[6748]=39779;
squeal_samples[6749]=35320;
squeal_samples[6750]=31144;
squeal_samples[6751]=27239;
squeal_samples[6752]=23585;
squeal_samples[6753]=20163;
squeal_samples[6754]=16964;
squeal_samples[6755]=13970;
squeal_samples[6756]=11176;
squeal_samples[6757]=8550;
squeal_samples[6758]=7690;
squeal_samples[6759]=10692;
squeal_samples[6760]=13749;
squeal_samples[6761]=16678;
squeal_samples[6762]=19471;
squeal_samples[6763]=22158;
squeal_samples[6764]=24714;
squeal_samples[6765]=27169;
squeal_samples[6766]=29503;
squeal_samples[6767]=31744;
squeal_samples[6768]=33883;
squeal_samples[6769]=35929;
squeal_samples[6770]=37876;
squeal_samples[6771]=39751;
squeal_samples[6772]=41530;
squeal_samples[6773]=43238;
squeal_samples[6774]=44863;
squeal_samples[6775]=46415;
squeal_samples[6776]=47905;
squeal_samples[6777]=49319;
squeal_samples[6778]=50681;
squeal_samples[6779]=51766;
squeal_samples[6780]=48324;
squeal_samples[6781]=43315;
squeal_samples[6782]=38625;
squeal_samples[6783]=34237;
squeal_samples[6784]=30133;
squeal_samples[6785]=26289;
squeal_samples[6786]=22701;
squeal_samples[6787]=19326;
squeal_samples[6788]=16188;
squeal_samples[6789]=13239;
squeal_samples[6790]=10488;
squeal_samples[6791]=7912;
squeal_samples[6792]=8308;
squeal_samples[6793]=11455;
squeal_samples[6794]=14483;
squeal_samples[6795]=17372;
squeal_samples[6796]=20146;
squeal_samples[6797]=22793;
squeal_samples[6798]=25328;
squeal_samples[6799]=27750;
squeal_samples[6800]=30063;
squeal_samples[6801]=32275;
squeal_samples[6802]=34391;
squeal_samples[6803]=36408;
squeal_samples[6804]=38347;
squeal_samples[6805]=40189;
squeal_samples[6806]=41954;
squeal_samples[6807]=43637;
squeal_samples[6808]=45244;
squeal_samples[6809]=46779;
squeal_samples[6810]=48250;
squeal_samples[6811]=49653;
squeal_samples[6812]=50996;
squeal_samples[6813]=51447;
squeal_samples[6814]=47029;
squeal_samples[6815]=42101;
squeal_samples[6816]=37487;
squeal_samples[6817]=33172;
squeal_samples[6818]=29128;
squeal_samples[6819]=25357;
squeal_samples[6820]=21819;
squeal_samples[6821]=18514;
squeal_samples[6822]=15417;
squeal_samples[6823]=12521;
squeal_samples[6824]=9817;
squeal_samples[6825]=7457;
squeal_samples[6826]=9095;
squeal_samples[6827]=12208;
squeal_samples[6828]=15204;
squeal_samples[6829]=18058;
squeal_samples[6830]=20807;
squeal_samples[6831]=23425;
squeal_samples[6832]=25928;
squeal_samples[6833]=28326;
squeal_samples[6834]=30604;
squeal_samples[6835]=32804;
squeal_samples[6836]=34889;
squeal_samples[6837]=36887;
squeal_samples[6838]=38799;
squeal_samples[6839]=40620;
squeal_samples[6840]=42365;
squeal_samples[6841]=44031;
squeal_samples[6842]=45621;
squeal_samples[6843]=47143;
squeal_samples[6844]=48592;
squeal_samples[6845]=49980;
squeal_samples[6846]=51308;
squeal_samples[6847]=50722;
squeal_samples[6848]=45757;
squeal_samples[6849]=40900;
squeal_samples[6850]=36370;
squeal_samples[6851]=32123;
squeal_samples[6852]=28151;
squeal_samples[6853]=24436;
squeal_samples[6854]=20959;
squeal_samples[6855]=17706;
squeal_samples[6856]=14662;
squeal_samples[6857]=11810;
squeal_samples[6858]=9158;
squeal_samples[6859]=7369;
squeal_samples[6860]=9871;
squeal_samples[6861]=12962;
squeal_samples[6862]=15912;
squeal_samples[6863]=18751;
squeal_samples[6864]=21458;
squeal_samples[6865]=24048;
squeal_samples[6866]=26526;
squeal_samples[6867]=28887;
squeal_samples[6868]=31158;
squeal_samples[6869]=33315;
squeal_samples[6870]=35391;
squeal_samples[6871]=37361;
squeal_samples[6872]=39252;
squeal_samples[6873]=41053;
squeal_samples[6874]=42775;
squeal_samples[6875]=44424;
squeal_samples[6876]=45994;
squeal_samples[6877]=47500;
squeal_samples[6878]=48931;
squeal_samples[6879]=50305;
squeal_samples[6880]=51614;
squeal_samples[6881]=49593;
squeal_samples[6882]=44496;
squeal_samples[6883]=39727;
squeal_samples[6884]=35268;
squeal_samples[6885]=31090;
squeal_samples[6886]=27187;
squeal_samples[6887]=23533;
squeal_samples[6888]=20107;
squeal_samples[6889]=16916;
squeal_samples[6890]=13915;
squeal_samples[6891]=11123;
squeal_samples[6892]=8498;
squeal_samples[6893]=7635;
squeal_samples[6894]=10643;
squeal_samples[6895]=13694;
squeal_samples[6896]=16626;
squeal_samples[6897]=19417;
squeal_samples[6898]=22106;
squeal_samples[6899]=24662;
squeal_samples[6900]=27115;
squeal_samples[6901]=29452;
squeal_samples[6902]=31688;
squeal_samples[6903]=33834;
squeal_samples[6904]=35873;
squeal_samples[6905]=37826;
squeal_samples[6906]=39696;
squeal_samples[6907]=41478;
squeal_samples[6908]=43186;
squeal_samples[6909]=44808;
squeal_samples[6910]=46364;
squeal_samples[6911]=47852;
squeal_samples[6912]=49265;
squeal_samples[6913]=50631;
squeal_samples[6914]=51709;
squeal_samples[6915]=48275;
squeal_samples[6916]=43260;
squeal_samples[6917]=38572;
squeal_samples[6918]=34187;
squeal_samples[6919]=30076;
squeal_samples[6920]=26240;
squeal_samples[6921]=22645;
squeal_samples[6922]=19274;
squeal_samples[6923]=16136;
squeal_samples[6924]=13185;
squeal_samples[6925]=10437;
squeal_samples[6926]=7857;
squeal_samples[6927]=8255;
squeal_samples[6928]=11404;
squeal_samples[6929]=14428;
squeal_samples[6930]=17323;
squeal_samples[6931]=20088;
squeal_samples[6932]=22744;
squeal_samples[6933]=25273;
squeal_samples[6934]=27700;
squeal_samples[6935]=30007;
squeal_samples[6936]=32225;
squeal_samples[6937]=34334;
squeal_samples[6938]=36360;
squeal_samples[6939]=38290;
squeal_samples[6940]=40139;
squeal_samples[6941]=41898;
squeal_samples[6942]=43586;
squeal_samples[6943]=45190;
squeal_samples[6944]=46726;
squeal_samples[6945]=48198;
squeal_samples[6946]=49597;
squeal_samples[6947]=50945;
squeal_samples[6948]=51755;
squeal_samples[6949]=47768;
squeal_samples[6950]=42783;
squeal_samples[6951]=38126;
squeal_samples[6952]=33764;
squeal_samples[6953]=29678;
squeal_samples[6954]=25869;
squeal_samples[6955]=22294;
squeal_samples[6956]=18952;
squeal_samples[6957]=15828;
squeal_samples[6958]=12902;
squeal_samples[6959]=10164;
squeal_samples[6960]=7653;
squeal_samples[6961]=8706;
squeal_samples[6962]=11843;
squeal_samples[6963]=14843;
squeal_samples[6964]=17721;
squeal_samples[6965]=20468;
squeal_samples[6966]=23104;
squeal_samples[6967]=25618;
squeal_samples[6968]=28029;
squeal_samples[6969]=30317;
squeal_samples[6970]=32530;
squeal_samples[6971]=34621;
squeal_samples[6972]=36637;
squeal_samples[6973]=38548;
squeal_samples[6974]=40383;
squeal_samples[6975]=42140;
squeal_samples[6976]=43805;
squeal_samples[6977]=45410;
squeal_samples[6978]=46928;
squeal_samples[6979]=48395;
squeal_samples[6980]=49783;
squeal_samples[6981]=51119;
squeal_samples[6982]=51565;
squeal_samples[6983]=47133;
squeal_samples[6984]=42189;
squeal_samples[6985]=37571;
squeal_samples[6986]=33242;
squeal_samples[6987]=29197;
squeal_samples[6988]=25411;
squeal_samples[6989]=21870;
squeal_samples[6990]=18549;
squeal_samples[6991]=15448;
squeal_samples[6992]=12549;
squeal_samples[6993]=9834;
squeal_samples[6994]=7476;
squeal_samples[6995]=9107;
squeal_samples[6996]=12220;
squeal_samples[6997]=15211;
squeal_samples[6998]=18064;
squeal_samples[6999]=20806;
squeal_samples[7000]=23417;
squeal_samples[7001]=25925;
squeal_samples[7002]=28308;
squeal_samples[7003]=30603;
squeal_samples[7004]=32783;
squeal_samples[7005]=34873;
squeal_samples[7006]=36869;
squeal_samples[7007]=38781;
squeal_samples[7008]=40598;
squeal_samples[7009]=42342;
squeal_samples[7010]=44002;
squeal_samples[7011]=45593;
squeal_samples[7012]=47114;
squeal_samples[7013]=48557;
squeal_samples[7014]=49949;
squeal_samples[7015]=51270;
squeal_samples[7016]=51251;
squeal_samples[7017]=46486;
squeal_samples[7018]=41592;
squeal_samples[7019]=37007;
squeal_samples[7020]=32716;
squeal_samples[7021]=28696;
squeal_samples[7022]=24946;
squeal_samples[7023]=21430;
squeal_samples[7024]=18142;
squeal_samples[7025]=15064;
squeal_samples[7026]=12187;
squeal_samples[7027]=9498;
squeal_samples[7028]=7377;
squeal_samples[7029]=9494;
squeal_samples[7030]=12586;
squeal_samples[7031]=15561;
squeal_samples[7032]=18407;
squeal_samples[7033]=21125;
squeal_samples[7034]=23728;
squeal_samples[7035]=26219;
squeal_samples[7036]=28590;
squeal_samples[7037]=30865;
squeal_samples[7038]=33041;
squeal_samples[7039]=35115;
squeal_samples[7040]=37102;
squeal_samples[7041]=38999;
squeal_samples[7042]=40810;
squeal_samples[7043]=42537;
squeal_samples[7044]=44196;
squeal_samples[7045]=45776;
squeal_samples[7046]=47285;
squeal_samples[7047]=48725;
squeal_samples[7048]=50107;
squeal_samples[7049]=51422;
squeal_samples[7050]=50829;
squeal_samples[7051]=45844;
squeal_samples[7052]=40985;
squeal_samples[7053]=36441;
squeal_samples[7054]=32186;
squeal_samples[7055]=28201;
squeal_samples[7056]=24480;
squeal_samples[7057]=20995;
squeal_samples[7058]=17731;
squeal_samples[7059]=14682;
squeal_samples[7060]=11833;
squeal_samples[7061]=9160;
squeal_samples[7062]=7373;
squeal_samples[7063]=9876;
squeal_samples[7064]=12953;
squeal_samples[7065]=15914;
squeal_samples[7066]=18731;
squeal_samples[7067]=21449;
squeal_samples[7068]=24029;
squeal_samples[7069]=26515;
squeal_samples[7070]=28866;
squeal_samples[7071]=31132;
squeal_samples[7072]=33292;
squeal_samples[7073]=35358;
squeal_samples[7074]=37331;
squeal_samples[7075]=39216;
squeal_samples[7076]=41017;
squeal_samples[7077]=42738;
squeal_samples[7078]=44384;
squeal_samples[7079]=45951;
squeal_samples[7080]=47457;
squeal_samples[7081]=48886;
squeal_samples[7082]=50256;
squeal_samples[7083]=51569;
squeal_samples[7084]=50303;
squeal_samples[7085]=45206;
squeal_samples[7086]=40386;
squeal_samples[7087]=35879;
squeal_samples[7088]=31656;
squeal_samples[7089]=27716;
squeal_samples[7090]=24016;
squeal_samples[7091]=20563;
squeal_samples[7092]=17328;
squeal_samples[7093]=14299;
squeal_samples[7094]=11476;
squeal_samples[7095]=8828;
squeal_samples[7096]=7452;
squeal_samples[7097]=10251;
squeal_samples[7098]=13321;
squeal_samples[7099]=16252;
squeal_samples[7100]=19072;
squeal_samples[7101]=21760;
squeal_samples[7102]=24338;
squeal_samples[7103]=26794;
squeal_samples[7104]=29146;
squeal_samples[7105]=31391;
squeal_samples[7106]=33542;
squeal_samples[7107]=35598;
squeal_samples[7108]=37558;
squeal_samples[7109]=39435;
squeal_samples[7110]=41228;
squeal_samples[7111]=42936;
squeal_samples[7112]=44571;
squeal_samples[7113]=46134;
squeal_samples[7114]=47622;
squeal_samples[7115]=49054;
squeal_samples[7116]=50410;
squeal_samples[7117]=51714;
squeal_samples[7118]=49682;
squeal_samples[7119]=44572;
squeal_samples[7120]=39799;
squeal_samples[7121]=35319;
squeal_samples[7122]=31141;
squeal_samples[7123]=27222;
squeal_samples[7124]=23561;
squeal_samples[7125]=20130;
squeal_samples[7126]=16923;
squeal_samples[7127]=13922;
squeal_samples[7128]=11121;
squeal_samples[7129]=8494;
squeal_samples[7130]=7624;
squeal_samples[7131]=10630;
squeal_samples[7132]=13679;
squeal_samples[7133]=16602;
squeal_samples[7134]=19398;
squeal_samples[7135]=22075;
squeal_samples[7136]=24637;
squeal_samples[7137]=27081;
squeal_samples[7138]=29413;
squeal_samples[7139]=31659;
squeal_samples[7140]=33784;
squeal_samples[7141]=35840;
squeal_samples[7142]=37779;
squeal_samples[7143]=39653;
squeal_samples[7144]=41430;
squeal_samples[7145]=43129;
squeal_samples[7146]=44761;
squeal_samples[7147]=46308;
squeal_samples[7148]=47798;
squeal_samples[7149]=49209;
squeal_samples[7150]=50570;
squeal_samples[7151]=51809;
squeal_samples[7152]=49010;
squeal_samples[7153]=43947;
squeal_samples[7154]=39207;
squeal_samples[7155]=34770;
squeal_samples[7156]=30624;
squeal_samples[7157]=26740;
squeal_samples[7158]=23109;
squeal_samples[7159]=19703;
squeal_samples[7160]=16524;
squeal_samples[7161]=13553;
squeal_samples[7162]=10769;
squeal_samples[7163]=8166;
squeal_samples[7164]=7881;
squeal_samples[7165]=11005;
squeal_samples[7166]=14039;
squeal_samples[7167]=16950;
squeal_samples[7168]=19723;
squeal_samples[7169]=22391;
squeal_samples[7170]=24931;
squeal_samples[7171]=27368;
squeal_samples[7172]=29688;
squeal_samples[7173]=31914;
squeal_samples[7174]=34036;
squeal_samples[7175]=36066;
squeal_samples[7176]=38009;
squeal_samples[7177]=39861;
squeal_samples[7178]=41632;
squeal_samples[7179]=43327;
squeal_samples[7180]=44936;
squeal_samples[7181]=46487;
squeal_samples[7182]=47959;
squeal_samples[7183]=49367;
squeal_samples[7184]=50720;
squeal_samples[7185]=51794;
squeal_samples[7186]=48348;
squeal_samples[7187]=43323;
squeal_samples[7188]=38624;
squeal_samples[7189]=34226;
squeal_samples[7190]=30108;
squeal_samples[7191]=26258;
squeal_samples[7192]=22659;
squeal_samples[7193]=19283;
squeal_samples[7194]=16133;
squeal_samples[7195]=13176;
squeal_samples[7196]=10425;
squeal_samples[7197]=7837;
squeal_samples[7198]=8232;
squeal_samples[7199]=11374;
squeal_samples[7200]=14398;
squeal_samples[7201]=17287;
squeal_samples[7202]=20050;
squeal_samples[7203]=22701;
squeal_samples[7204]=25229;
squeal_samples[7205]=27653;
squeal_samples[7206]=29956;
squeal_samples[7207]=32173;
squeal_samples[7208]=34284;
squeal_samples[7209]=36301;
squeal_samples[7210]=38232;
squeal_samples[7211]=40071;
squeal_samples[7212]=41842;
squeal_samples[7213]=43513;
squeal_samples[7214]=45127;
squeal_samples[7215]=46656;
squeal_samples[7216]=48129;
squeal_samples[7217]=49527;
squeal_samples[7218]=50869;
squeal_samples[7219]=51681;
squeal_samples[7220]=47685;
squeal_samples[7221]=42707;
squeal_samples[7222]=38048;
squeal_samples[7223]=33677;
squeal_samples[7224]=29605;
squeal_samples[7225]=25780;
squeal_samples[7226]=22213;
squeal_samples[7227]=18863;
squeal_samples[7228]=15737;
squeal_samples[7229]=12808;
squeal_samples[7230]=10076;
squeal_samples[7231]=7563;
squeal_samples[7232]=8616;
squeal_samples[7233]=11751;
squeal_samples[7234]=14749;
squeal_samples[7235]=17631;
squeal_samples[7236]=20377;
squeal_samples[7237]=23009;
squeal_samples[7238]=25526;
squeal_samples[7239]=27925;
squeal_samples[7240]=30227;
squeal_samples[7241]=32426;
squeal_samples[7242]=34524;
squeal_samples[7243]=36535;
squeal_samples[7244]=38454;
squeal_samples[7245]=40284;
squeal_samples[7246]=42039;
squeal_samples[7247]=43706;
squeal_samples[7248]=45308;
squeal_samples[7249]=46836;
squeal_samples[7250]=48293;
squeal_samples[7251]=49685;
squeal_samples[7252]=51017;
squeal_samples[7253]=51467;
squeal_samples[7254]=47031;
squeal_samples[7255]=42092;
squeal_samples[7256]=37468;
squeal_samples[7257]=33145;
squeal_samples[7258]=29095;
squeal_samples[7259]=25307;
squeal_samples[7260]=21770;
squeal_samples[7261]=18448;
squeal_samples[7262]=15350;
squeal_samples[7263]=12446;
squeal_samples[7264]=9738;
squeal_samples[7265]=7372;
squeal_samples[7266]=9005;
squeal_samples[7267]=12113;
squeal_samples[7268]=15106;
squeal_samples[7269]=17959;
squeal_samples[7270]=20699;
squeal_samples[7271]=23314;
squeal_samples[7272]=25817;
squeal_samples[7273]=28207;
squeal_samples[7274]=30492;
squeal_samples[7275]=32689;
squeal_samples[7276]=34767;
squeal_samples[7277]=36769;
squeal_samples[7278]=38673;
squeal_samples[7279]=40498;
squeal_samples[7280]=42238;
squeal_samples[7281]=43899;
squeal_samples[7282]=45490;
squeal_samples[7283]=47008;
squeal_samples[7284]=48457;
squeal_samples[7285]=49847;
squeal_samples[7286]=51165;
squeal_samples[7287]=51607;
squeal_samples[7288]=47164;
squeal_samples[7289]=42213;
squeal_samples[7290]=37586;
squeal_samples[7291]=33246;
squeal_samples[7292]=29189;
squeal_samples[7293]=25398;
squeal_samples[7294]=21847;
squeal_samples[7295]=18529;
squeal_samples[7296]=15417;
squeal_samples[7297]=12510;
squeal_samples[7298]=9793;
squeal_samples[7299]=7427;
squeal_samples[7300]=9053;
squeal_samples[7301]=12169;
squeal_samples[7302]=15148;
squeal_samples[7303]=18010;
squeal_samples[7304]=20742;
squeal_samples[7305]=23357;
squeal_samples[7306]=25858;
squeal_samples[7307]=28239;
squeal_samples[7308]=30530;
squeal_samples[7309]=32709;
squeal_samples[7310]=34801;
squeal_samples[7311]=36793;
squeal_samples[7312]=38700;
squeal_samples[7313]=40519;
squeal_samples[7314]=42259;
squeal_samples[7315]=43923;
squeal_samples[7316]=45505;
squeal_samples[7317]=47024;
squeal_samples[7318]=48471;
squeal_samples[7319]=49860;
squeal_samples[7320]=51181;
squeal_samples[7321]=51619;
squeal_samples[7322]=47173;
squeal_samples[7323]=42222;
squeal_samples[7324]=37588;
squeal_samples[7325]=33257;
squeal_samples[7326]=29194;
squeal_samples[7327]=25411;
squeal_samples[7328]=21846;
squeal_samples[7329]=18530;
squeal_samples[7330]=15418;
squeal_samples[7331]=12514;
squeal_samples[7332]=9796;
squeal_samples[7333]=7430;
squeal_samples[7334]=9051;
squeal_samples[7335]=12166;
squeal_samples[7336]=15148;
squeal_samples[7337]=18005;
squeal_samples[7338]=20736;
squeal_samples[7339]=23354;
squeal_samples[7340]=25850;
squeal_samples[7341]=28238;
squeal_samples[7342]=30526;
squeal_samples[7343]=32703;
squeal_samples[7344]=34797;
squeal_samples[7345]=36787;
squeal_samples[7346]=38691;
squeal_samples[7347]=40517;
squeal_samples[7348]=42251;
squeal_samples[7349]=43914;
squeal_samples[7350]=45501;
squeal_samples[7351]=47012;
squeal_samples[7352]=48467;
squeal_samples[7353]=49848;
squeal_samples[7354]=51176;
squeal_samples[7355]=51610;
squeal_samples[7356]=47167;
squeal_samples[7357]=42212;
squeal_samples[7358]=37583;
squeal_samples[7359]=33245;
squeal_samples[7360]=29185;
squeal_samples[7361]=25395;
squeal_samples[7362]=21841;
squeal_samples[7363]=18519;
squeal_samples[7364]=15407;
squeal_samples[7365]=12500;
squeal_samples[7366]=9784;
squeal_samples[7367]=7416;
squeal_samples[7368]=9038;
squeal_samples[7369]=12152;
squeal_samples[7370]=15136;
squeal_samples[7371]=17991;
squeal_samples[7372]=20730;
squeal_samples[7373]=23338;
squeal_samples[7374]=25845;
squeal_samples[7375]=28224;
squeal_samples[7376]=30511;
squeal_samples[7377]=32694;
squeal_samples[7378]=34780;
squeal_samples[7379]=36776;
squeal_samples[7380]=38677;
squeal_samples[7381]=40504;
squeal_samples[7382]=42239;
squeal_samples[7383]=43900;
squeal_samples[7384]=45488;
squeal_samples[7385]=47005;
squeal_samples[7386]=48452;
squeal_samples[7387]=49839;
squeal_samples[7388]=51158;
squeal_samples[7389]=51602;
squeal_samples[7390]=47148;
squeal_samples[7391]=42205;
squeal_samples[7392]=37564;
squeal_samples[7393]=33239;
squeal_samples[7394]=29172;
squeal_samples[7395]=25384;
squeal_samples[7396]=21827;
squeal_samples[7397]=18507;
squeal_samples[7398]=15394;
squeal_samples[7399]=12487;
squeal_samples[7400]=9770;
squeal_samples[7401]=7404;
squeal_samples[7402]=9029;
squeal_samples[7403]=12141;
squeal_samples[7404]=15120;
squeal_samples[7405]=17981;
squeal_samples[7406]=20714;
squeal_samples[7407]=23328;
squeal_samples[7408]=25829;
squeal_samples[7409]=28212;
squeal_samples[7410]=30499;
squeal_samples[7411]=32678;
squeal_samples[7412]=34770;
squeal_samples[7413]=36761;
squeal_samples[7414]=38665;
squeal_samples[7415]=40491;
squeal_samples[7416]=42224;
squeal_samples[7417]=43890;
squeal_samples[7418]=45472;
squeal_samples[7419]=46993;
squeal_samples[7420]=48441;
squeal_samples[7421]=49822;
squeal_samples[7422]=51149;
squeal_samples[7423]=51585;
squeal_samples[7424]=47138;
squeal_samples[7425]=42191;
squeal_samples[7426]=37551;
squeal_samples[7427]=33224;
squeal_samples[7428]=29160;
squeal_samples[7429]=25372;
squeal_samples[7430]=21813;
squeal_samples[7431]=18495;
squeal_samples[7432]=15383;
squeal_samples[7433]=12477;
squeal_samples[7434]=9755;
squeal_samples[7435]=7392;
squeal_samples[7436]=9017;
squeal_samples[7437]=12125;
squeal_samples[7438]=15111;
squeal_samples[7439]=17964;
squeal_samples[7440]=20704;
squeal_samples[7441]=23312;
squeal_samples[7442]=25820;
squeal_samples[7443]=28196;
squeal_samples[7444]=30487;
squeal_samples[7445]=32666;
squeal_samples[7446]=34755;
squeal_samples[7447]=36749;
squeal_samples[7448]=38653;
squeal_samples[7449]=40474;
squeal_samples[7450]=42218;
squeal_samples[7451]=43869;
squeal_samples[7452]=45465;
squeal_samples[7453]=46977;
squeal_samples[7454]=48427;
squeal_samples[7455]=49812;
squeal_samples[7456]=51133;
squeal_samples[7457]=51574;
squeal_samples[7458]=47124;
squeal_samples[7459]=42177;
squeal_samples[7460]=37540;
squeal_samples[7461]=33209;
squeal_samples[7462]=29149;
squeal_samples[7463]=25356;
squeal_samples[7464]=21803;
squeal_samples[7465]=18479;
squeal_samples[7466]=15374;
squeal_samples[7467]=12460;
squeal_samples[7468]=9744;
squeal_samples[7469]=7379;
squeal_samples[7470]=9003;
squeal_samples[7471]=12114;
squeal_samples[7472]=15095;
squeal_samples[7473]=17953;
squeal_samples[7474]=20689;
squeal_samples[7475]=23303;
squeal_samples[7476]=25801;
squeal_samples[7477]=28189;
squeal_samples[7478]=30469;
squeal_samples[7479]=32655;
squeal_samples[7480]=34743;
squeal_samples[7481]=36733;
squeal_samples[7482]=38642;
squeal_samples[7483]=40462;
squeal_samples[7484]=42201;
squeal_samples[7485]=43861;
squeal_samples[7486]=45448;
squeal_samples[7487]=46966;
squeal_samples[7488]=48414;
squeal_samples[7489]=49797;
squeal_samples[7490]=51123;
squeal_samples[7491]=51558;
squeal_samples[7492]=47116;
squeal_samples[7493]=42157;
squeal_samples[7494]=37534;
squeal_samples[7495]=33189;
squeal_samples[7496]=29143;
squeal_samples[7497]=25338;
squeal_samples[7498]=21792;
squeal_samples[7499]=18466;
squeal_samples[7500]=15359;
squeal_samples[7501]=12449;
squeal_samples[7502]=9731;
squeal_samples[7503]=7364;
squeal_samples[7504]=8992;
squeal_samples[7505]=12100;
squeal_samples[7506]=15081;
squeal_samples[7507]=17944;
squeal_samples[7508]=20671;
squeal_samples[7509]=23293;
squeal_samples[7510]=25788;
squeal_samples[7511]=28174;
squeal_samples[7512]=30458;
squeal_samples[7513]=32642;
squeal_samples[7514]=34728;
squeal_samples[7515]=36724;
squeal_samples[7516]=38625;
squeal_samples[7517]=40451;
squeal_samples[7518]=42187;
squeal_samples[7519]=43850;
squeal_samples[7520]=45432;
squeal_samples[7521]=46956;
squeal_samples[7522]=48398;
squeal_samples[7523]=49787;
squeal_samples[7524]=51108;
squeal_samples[7525]=51546;
squeal_samples[7526]=47100;
squeal_samples[7527]=42149;
squeal_samples[7528]=37515;
squeal_samples[7529]=33183;
squeal_samples[7530]=29124;
squeal_samples[7531]=25328;
squeal_samples[7532]=21779;
squeal_samples[7533]=18451;
squeal_samples[7534]=15349;
squeal_samples[7535]=12434;
squeal_samples[7536]=9719;
squeal_samples[7537]=7350;
squeal_samples[7538]=8980;
squeal_samples[7539]=12086;
squeal_samples[7540]=15069;
squeal_samples[7541]=17930;
squeal_samples[7542]=20659;
squeal_samples[7543]=23279;
squeal_samples[7544]=25775;
squeal_samples[7545]=28161;
squeal_samples[7546]=30447;
squeal_samples[7547]=32625;
squeal_samples[7548]=34719;
squeal_samples[7549]=36707;
squeal_samples[7550]=38616;
squeal_samples[7551]=40435;
squeal_samples[7552]=42176;
squeal_samples[7553]=43835;
squeal_samples[7554]=45421;
squeal_samples[7555]=46942;
squeal_samples[7556]=48385;
squeal_samples[7557]=49774;
squeal_samples[7558]=51095;
squeal_samples[7559]=51534;
squeal_samples[7560]=47086;
squeal_samples[7561]=42137;
squeal_samples[7562]=37501;
squeal_samples[7563]=33171;
squeal_samples[7564]=29109;
squeal_samples[7565]=25318;
squeal_samples[7566]=21763;
squeal_samples[7567]=18441;
squeal_samples[7568]=15334;
squeal_samples[7569]=12421;
squeal_samples[7570]=9707;
squeal_samples[7571]=7337;
squeal_samples[7572]=8967;
squeal_samples[7573]=12071;
squeal_samples[7574]=15061;
squeal_samples[7575]=17910;
squeal_samples[7576]=20653;
squeal_samples[7577]=23261;
squeal_samples[7578]=25764;
squeal_samples[7579]=28149;
squeal_samples[7580]=30431;
squeal_samples[7581]=32615;
squeal_samples[7582]=34704;
squeal_samples[7583]=36696;
squeal_samples[7584]=38600;
squeal_samples[7585]=40425;
squeal_samples[7586]=42160;
squeal_samples[7587]=43825;
squeal_samples[7588]=45405;
squeal_samples[7589]=46932;
squeal_samples[7590]=48370;
squeal_samples[7591]=49763;
squeal_samples[7592]=51080;
squeal_samples[7593]=51522;
squeal_samples[7594]=47072;
squeal_samples[7595]=42125;
squeal_samples[7596]=37488;
squeal_samples[7597]=33157;
squeal_samples[7598]=29098;
squeal_samples[7599]=25303;
squeal_samples[7600]=21750;
squeal_samples[7601]=18428;
squeal_samples[7602]=15321;
squeal_samples[7603]=12409;
squeal_samples[7604]=9692;
squeal_samples[7605]=7326;
squeal_samples[7606]=8951;
squeal_samples[7607]=12062;
squeal_samples[7608]=15043;
squeal_samples[7609]=17902;
squeal_samples[7610]=20636;
squeal_samples[7611]=23251;
squeal_samples[7612]=25748;
squeal_samples[7613]=28138;
squeal_samples[7614]=30416;
squeal_samples[7615]=32604;
squeal_samples[7616]=34690;
squeal_samples[7617]=36682;
squeal_samples[7618]=38589;
squeal_samples[7619]=40409;
squeal_samples[7620]=42151;
squeal_samples[7621]=43807;
squeal_samples[7622]=45397;
squeal_samples[7623]=46913;
squeal_samples[7624]=48363;
squeal_samples[7625]=49743;
squeal_samples[7626]=51072;
squeal_samples[7627]=51862;
squeal_samples[7628]=47851;
squeal_samples[7629]=42848;
squeal_samples[7630]=38167;
squeal_samples[7631]=33787;
squeal_samples[7632]=29690;
squeal_samples[7633]=25853;
squeal_samples[7634]=22265;
squeal_samples[7635]=18909;
squeal_samples[7636]=15768;
squeal_samples[7637]=12832;
squeal_samples[7638]=10080;
squeal_samples[7639]=7558;
squeal_samples[7640]=8600;
squeal_samples[7641]=11735;
squeal_samples[7642]=14723;
squeal_samples[7643]=17598;
squeal_samples[7644]=20340;
squeal_samples[7645]=22970;
squeal_samples[7646]=25483;
squeal_samples[7647]=27878;
squeal_samples[7648]=30171;
squeal_samples[7649]=32369;
squeal_samples[7650]=34462;
squeal_samples[7651]=36472;
squeal_samples[7652]=38383;
squeal_samples[7653]=40215;
squeal_samples[7654]=41954;
squeal_samples[7655]=43630;
squeal_samples[7656]=45222;
squeal_samples[7657]=46747;
squeal_samples[7658]=48199;
squeal_samples[7659]=49592;
squeal_samples[7660]=50919;
squeal_samples[7661]=51983;
squeal_samples[7662]=48509;
squeal_samples[7663]=43467;
squeal_samples[7664]=38744;
squeal_samples[7665]=34325;
squeal_samples[7666]=30191;
squeal_samples[7667]=26323;
squeal_samples[7668]=22710;
squeal_samples[7669]=19316;
squeal_samples[7670]=16150;
squeal_samples[7671]=13187;
squeal_samples[7672]=10413;
squeal_samples[7673]=7825;
squeal_samples[7674]=8200;
squeal_samples[7675]=11344;
squeal_samples[7676]=14359;
squeal_samples[7677]=17234;
squeal_samples[7678]=20008;
squeal_samples[7679]=22638;
squeal_samples[7680]=25175;
squeal_samples[7681]=27578;
squeal_samples[7682]=29893;
squeal_samples[7683]=32089;
squeal_samples[7684]=34204;
squeal_samples[7685]=36219;
squeal_samples[7686]=38141;
squeal_samples[7687]=39980;
squeal_samples[7688]=41736;
squeal_samples[7689]=43413;
squeal_samples[7690]=45023;
squeal_samples[7691]=46551;
squeal_samples[7692]=48015;
squeal_samples[7693]=49409;
squeal_samples[7694]=50749;
squeal_samples[7695]=51974;
squeal_samples[7696]=49155;
squeal_samples[7697]=44066;
squeal_samples[7698]=39311;
squeal_samples[7699]=34849;
squeal_samples[7700]=30689;
squeal_samples[7701]=26779;
squeal_samples[7702]=23138;
squeal_samples[7703]=19718;
squeal_samples[7704]=16525;
squeal_samples[7705]=13538;
squeal_samples[7706]=10740;
squeal_samples[7707]=8130;
squeal_samples[7708]=7829;
squeal_samples[7709]=10948;
squeal_samples[7710]=13975;
squeal_samples[7711]=16882;
squeal_samples[7712]=19650;
squeal_samples[7713]=22312;
squeal_samples[7714]=24846;
squeal_samples[7715]=27277;
squeal_samples[7716]=29594;
squeal_samples[7717]=31812;
squeal_samples[7718]=33931;
squeal_samples[7719]=35960;
squeal_samples[7720]=37889;
squeal_samples[7721]=39746;
squeal_samples[7722]=41510;
squeal_samples[7723]=43201;
squeal_samples[7724]=44813;
squeal_samples[7725]=46349;
squeal_samples[7726]=47821;
squeal_samples[7727]=49229;
squeal_samples[7728]=50573;
squeal_samples[7729]=51856;
squeal_samples[7730]=49808;
squeal_samples[7731]=44670;
squeal_samples[7732]=39873;
squeal_samples[7733]=35379;
squeal_samples[7734]=31173;
squeal_samples[7735]=27252;
squeal_samples[7736]=23564;
squeal_samples[7737]=20122;
squeal_samples[7738]=16895;
squeal_samples[7739]=13886;
squeal_samples[7740]=11067;
squeal_samples[7741]=8433;
squeal_samples[7742]=7552;
squeal_samples[7743]=10545;
squeal_samples[7744]=13593;
squeal_samples[7745]=16504;
squeal_samples[7746]=19300;
squeal_samples[7747]=21971;
squeal_samples[7748]=24519;
squeal_samples[7749]=26967;
squeal_samples[7750]=29290;
squeal_samples[7751]=31531;
squeal_samples[7752]=33655;
squeal_samples[7753]=35698;
squeal_samples[7754]=37646;
squeal_samples[7755]=39500;
squeal_samples[7756]=41284;
squeal_samples[7757]=42973;
squeal_samples[7758]=44602;
squeal_samples[7759]=46149;
squeal_samples[7760]=47631;
squeal_samples[7761]=49040;
squeal_samples[7762]=50397;
squeal_samples[7763]=51688;
squeal_samples[7764]=50398;
squeal_samples[7765]=45288;
squeal_samples[7766]=40443;
squeal_samples[7767]=35915;
squeal_samples[7768]=31674;
squeal_samples[7769]=27707;
squeal_samples[7770]=24000;
squeal_samples[7771]=20524;
squeal_samples[7772]=17276;
squeal_samples[7773]=14240;
squeal_samples[7774]=11399;
squeal_samples[7775]=8741;
squeal_samples[7776]=7350;
squeal_samples[7777]=10147;
squeal_samples[7778]=13203;
squeal_samples[7779]=16140;
squeal_samples[7780]=18942;
squeal_samples[7781]=21631;
squeal_samples[7782]=24200;
squeal_samples[7783]=26650;
squeal_samples[7784]=29001;
squeal_samples[7785]=31238;
squeal_samples[7786]=33383;
squeal_samples[7787]=35436;
squeal_samples[7788]=37391;
squeal_samples[7789]=39263;
squeal_samples[7790]=41051;
squeal_samples[7791]=42757;
squeal_samples[7792]=44390;
squeal_samples[7793]=45950;
squeal_samples[7794]=47434;
squeal_samples[7795]=48859;
squeal_samples[7796]=50210;
squeal_samples[7797]=51519;
squeal_samples[7798]=50902;
squeal_samples[7799]=45899;
squeal_samples[7800]=41018;
squeal_samples[7801]=36451;
squeal_samples[7802]=32174;
squeal_samples[7803]=28175;
squeal_samples[7804]=24436;
squeal_samples[7805]=20936;
squeal_samples[7806]=17659;
squeal_samples[7807]=14597;
squeal_samples[7808]=11727;
squeal_samples[7809]=9050;
squeal_samples[7810]=7246;
squeal_samples[7811]=9740;
squeal_samples[7812]=12818;
squeal_samples[7813]=15767;
squeal_samples[7814]=18586;
squeal_samples[7815]=21289;
squeal_samples[7816]=23870;
squeal_samples[7817]=26342;
squeal_samples[7818]=28698;
squeal_samples[7819]=30953;
squeal_samples[7820]=33111;
squeal_samples[7821]=35171;
squeal_samples[7822]=37138;
squeal_samples[7823]=39019;
squeal_samples[7824]=40817;
squeal_samples[7825]=42538;
squeal_samples[7826]=44175;
squeal_samples[7827]=45743;
squeal_samples[7828]=47236;
squeal_samples[7829]=48671;
squeal_samples[7830]=50037;
squeal_samples[7831]=51345;
squeal_samples[7832]=51299;
squeal_samples[7833]=46520;
squeal_samples[7834]=41598;
squeal_samples[7835]=36991;
squeal_samples[7836]=32679;
squeal_samples[7837]=28650;
squeal_samples[7838]=24879;
squeal_samples[7839]=21347;
squeal_samples[7840]=18041;
squeal_samples[7841]=14956;
squeal_samples[7842]=12061;
squeal_samples[7843]=9362;
squeal_samples[7844]=7229;
squeal_samples[7845]=9334;
squeal_samples[7846]=12428;
squeal_samples[7847]=15391;
squeal_samples[7848]=18230;
squeal_samples[7849]=20941;
squeal_samples[7850]=23546;
squeal_samples[7851]=26021;
squeal_samples[7852]=28395;
squeal_samples[7853]=30662;
squeal_samples[7854]=32833;
squeal_samples[7855]=34903;
squeal_samples[7856]=36885;
squeal_samples[7857]=38780;
squeal_samples[7858]=40586;
squeal_samples[7859]=42313;
squeal_samples[7860]=43963;
squeal_samples[7861]=45537;
squeal_samples[7862]=47043;
squeal_samples[7863]=48480;
squeal_samples[7864]=49858;
squeal_samples[7865]=51168;
squeal_samples[7866]=51601;
squeal_samples[7867]=47144;
squeal_samples[7868]=42182;
squeal_samples[7869]=37538;
squeal_samples[7870]=33193;
squeal_samples[7871]=29125;
squeal_samples[7872]=25324;
squeal_samples[7873]=21761;
squeal_samples[7874]=18433;
squeal_samples[7875]=15314;
squeal_samples[7876]=12404;
squeal_samples[7877]=9675;
squeal_samples[7878]=7303;
squeal_samples[7879]=8925;
squeal_samples[7880]=12033;
squeal_samples[7881]=15017;
squeal_samples[7882]=17866;
squeal_samples[7883]=20601;
squeal_samples[7884]=23208;
squeal_samples[7885]=25710;
squeal_samples[7886]=28090;
squeal_samples[7887]=30368;
squeal_samples[7888]=32555;
squeal_samples[7889]=34633;
squeal_samples[7890]=36631;
squeal_samples[7891]=38532;
squeal_samples[7892]=40350;
squeal_samples[7893]=42090;
squeal_samples[7894]=43746;
squeal_samples[7895]=45339;
squeal_samples[7896]=46841;
squeal_samples[7897]=48297;
squeal_samples[7898]=49674;
squeal_samples[7899]=50998;
squeal_samples[7900]=51795;
squeal_samples[7901]=47772;
squeal_samples[7902]=42772;
squeal_samples[7903]=38092;
squeal_samples[7904]=33704;
squeal_samples[7905]=29609;
squeal_samples[7906]=25770;
squeal_samples[7907]=22186;
squeal_samples[7908]=18818;
squeal_samples[7909]=15686;
squeal_samples[7910]=12740;
squeal_samples[7911]=9996;
squeal_samples[7912]=7469;
squeal_samples[7913]=8515;
squeal_samples[7914]=11640;
squeal_samples[7915]=14634;
squeal_samples[7916]=17507;
squeal_samples[7917]=20250;
squeal_samples[7918]=22877;
squeal_samples[7919]=25390;
squeal_samples[7920]=27785;
squeal_samples[7921]=30080;
squeal_samples[7922]=32274;
squeal_samples[7923]=34368;
squeal_samples[7924]=36371;
squeal_samples[7925]=38286;
squeal_samples[7926]=40115;
squeal_samples[7927]=41866;
squeal_samples[7928]=43527;
squeal_samples[7929]=45130;
squeal_samples[7930]=46643;
squeal_samples[7931]=48105;
squeal_samples[7932]=49492;
squeal_samples[7933]=50823;
squeal_samples[7934]=51884;
squeal_samples[7935]=48411;
squeal_samples[7936]=43370;
squeal_samples[7937]=38639;
squeal_samples[7938]=34230;
squeal_samples[7939]=30090;
squeal_samples[7940]=26229;
squeal_samples[7941]=22603;
squeal_samples[7942]=19216;
squeal_samples[7943]=16051;
squeal_samples[7944]=13082;
squeal_samples[7945]=10313;
squeal_samples[7946]=7724;
squeal_samples[7947]=8099;
squeal_samples[7948]=11241;
squeal_samples[7949]=14258;
squeal_samples[7950]=17140;
squeal_samples[7951]=19900;
squeal_samples[7952]=22546;
squeal_samples[7953]=25065;
squeal_samples[7954]=27487;
squeal_samples[7955]=29784;
squeal_samples[7956]=31988;
squeal_samples[7957]=34102;
squeal_samples[7958]=36112;
squeal_samples[7959]=38040;
squeal_samples[7960]=39882;
squeal_samples[7961]=41631;
squeal_samples[7962]=43313;
squeal_samples[7963]=44916;
squeal_samples[7964]=46449;
squeal_samples[7965]=47910;
squeal_samples[7966]=49307;
squeal_samples[7967]=50645;
squeal_samples[7968]=51924;
squeal_samples[7969]=49861;
squeal_samples[7970]=44719;
squeal_samples[7971]=39911;
squeal_samples[7972]=35412;
squeal_samples[7973]=31200;
squeal_samples[7974]=27261;
squeal_samples[7975]=23575;
squeal_samples[7976]=20126;
squeal_samples[7977]=16894;
squeal_samples[7978]=13874;
squeal_samples[7979]=11055;
squeal_samples[7980]=8413;
squeal_samples[7981]=7526;
squeal_samples[7982]=10521;
squeal_samples[7983]=13565;
squeal_samples[7984]=16476;
squeal_samples[7985]=19269;
squeal_samples[7986]=21932;
squeal_samples[7987]=24488;
squeal_samples[7988]=26919;
squeal_samples[7989]=29255;
squeal_samples[7990]=31479;
squeal_samples[7991]=33611;
squeal_samples[7992]=35645;
squeal_samples[7993]=37591;
squeal_samples[7994]=39452;
squeal_samples[7995]=41221;
squeal_samples[7996]=42926;
squeal_samples[7997]=44540;
squeal_samples[7998]=46088;
squeal_samples[7999]=47571;
squeal_samples[8000]=48985;
squeal_samples[8001]=50329;
squeal_samples[8002]=51627;
squeal_samples[8003]=50997;
squeal_samples[8004]=45986;
squeal_samples[8005]=41090;
squeal_samples[8006]=36516;
squeal_samples[8007]=32231;
squeal_samples[8008]=28224;
squeal_samples[8009]=24477;
squeal_samples[8010]=20966;
squeal_samples[8011]=17686;
squeal_samples[8012]=14610;
squeal_samples[8013]=11743;
squeal_samples[8014]=9059;
squeal_samples[8015]=7249;
squeal_samples[8016]=9739;
squeal_samples[8017]=12812;
squeal_samples[8018]=15758;
squeal_samples[8019]=18576;
squeal_samples[8020]=21275;
squeal_samples[8021]=23852;
squeal_samples[8022]=26320;
squeal_samples[8023]=28673;
squeal_samples[8024]=30927;
squeal_samples[8025]=33081;
squeal_samples[8026]=35141;
squeal_samples[8027]=37111;
squeal_samples[8028]=38983;
squeal_samples[8029]=40786;
squeal_samples[8030]=42494;
squeal_samples[8031]=44140;
squeal_samples[8032]=45698;
squeal_samples[8033]=47202;
squeal_samples[8034]=48622;
squeal_samples[8035]=49993;
squeal_samples[8036]=51295;
squeal_samples[8037]=51714;
squeal_samples[8038]=47249;
squeal_samples[8039]=42273;
squeal_samples[8040]=37623;
squeal_samples[8041]=33265;
squeal_samples[8042]=29195;
squeal_samples[8043]=25382;
squeal_samples[8044]=21811;
squeal_samples[8045]=18477;
squeal_samples[8046]=15352;
squeal_samples[8047]=12431;
squeal_samples[8048]=9699;
squeal_samples[8049]=7318;
squeal_samples[8050]=8938;
squeal_samples[8051]=12042;
squeal_samples[8052]=15026;
squeal_samples[8053]=17869;
squeal_samples[8054]=20604;
squeal_samples[8055]=23202;
squeal_samples[8056]=25704;
squeal_samples[8057]=28081;
squeal_samples[8058]=30358;
squeal_samples[8059]=32544;
squeal_samples[8060]=34623;
squeal_samples[8061]=36614;
squeal_samples[8062]=38511;
squeal_samples[8063]=40330;
squeal_samples[8064]=42067;
squeal_samples[8065]=43722;
squeal_samples[8066]=45308;
squeal_samples[8067]=46817;
squeal_samples[8068]=48264;
squeal_samples[8069]=49641;
squeal_samples[8070]=50966;
squeal_samples[8071]=52018;
squeal_samples[8072]=48532;
squeal_samples[8073]=43475;
squeal_samples[8074]=38742;
squeal_samples[8075]=34315;
squeal_samples[8076]=30173;
squeal_samples[8077]=26298;
squeal_samples[8078]=22673;
squeal_samples[8079]=19278;
squeal_samples[8080]=16101;
squeal_samples[8081]=13130;
squeal_samples[8082]=10352;
squeal_samples[8083]=7755;
squeal_samples[8084]=8127;
squeal_samples[8085]=11267;
squeal_samples[8086]=14275;
squeal_samples[8087]=17161;
squeal_samples[8088]=19913;
squeal_samples[8089]=22552;
squeal_samples[8090]=25076;
squeal_samples[8091]=27487;
squeal_samples[8092]=29787;
squeal_samples[8093]=31993;
squeal_samples[8094]=34095;
squeal_samples[8095]=36114;
squeal_samples[8096]=38029;
squeal_samples[8097]=39874;
squeal_samples[8098]=41624;
squeal_samples[8099]=43302;
squeal_samples[8100]=44906;
squeal_samples[8101]=46434;
squeal_samples[8102]=47896;
squeal_samples[8103]=49294;
squeal_samples[8104]=50625;
squeal_samples[8105]=51900;
squeal_samples[8106]=49837;
squeal_samples[8107]=44694;
squeal_samples[8108]=39886;
squeal_samples[8109]=35386;
squeal_samples[8110]=31165;
squeal_samples[8111]=27235;
squeal_samples[8112]=23542;
squeal_samples[8113]=20093;
squeal_samples[8114]=16858;
squeal_samples[8115]=13841;
squeal_samples[8116]=11011;
squeal_samples[8117]=8380;
squeal_samples[8118]=7489;
squeal_samples[8119]=10481;
squeal_samples[8120]=13526;
squeal_samples[8121]=16433;
squeal_samples[8122]=19230;
squeal_samples[8123]=21891;
squeal_samples[8124]=24446;
squeal_samples[8125]=26881;
squeal_samples[8126]=29211;
squeal_samples[8127]=31437;
squeal_samples[8128]=33567;
squeal_samples[8129]=35605;
squeal_samples[8130]=37547;
squeal_samples[8131]=39409;
squeal_samples[8132]=41183;
squeal_samples[8133]=42878;
squeal_samples[8134]=44494;
squeal_samples[8135]=46042;
squeal_samples[8136]=47526;
squeal_samples[8137]=48937;
squeal_samples[8138]=50287;
squeal_samples[8139]=51576;
squeal_samples[8140]=50955;
squeal_samples[8141]=45936;
squeal_samples[8142]=41048;
squeal_samples[8143]=36467;
squeal_samples[8144]=32183;
squeal_samples[8145]=28174;
squeal_samples[8146]=24429;
squeal_samples[8147]=20919;
squeal_samples[8148]=17635;
squeal_samples[8149]=14564;
squeal_samples[8150]=11692;
squeal_samples[8151]=9005;
squeal_samples[8152]=7202;
squeal_samples[8153]=9689;
squeal_samples[8154]=12763;
squeal_samples[8155]=15705;
squeal_samples[8156]=18525;
squeal_samples[8157]=21223;
squeal_samples[8158]=23803;
squeal_samples[8159]=26271;
squeal_samples[8160]=28623;
squeal_samples[8161]=30879;
squeal_samples[8162]=33031;
squeal_samples[8163]=35092;
squeal_samples[8164]=37056;
squeal_samples[8165]=38935;
squeal_samples[8166]=40730;
squeal_samples[8167]=42447;
squeal_samples[8168]=44085;
squeal_samples[8169]=45651;
squeal_samples[8170]=47146;
squeal_samples[8171]=48579;
squeal_samples[8172]=49941;
squeal_samples[8173]=51247;
squeal_samples[8174]=51665;
squeal_samples[8175]=47195;
squeal_samples[8176]=42225;
squeal_samples[8177]=37572;
squeal_samples[8178]=33221;
squeal_samples[8179]=29136;
squeal_samples[8180]=25335;
squeal_samples[8181]=21758;
squeal_samples[8182]=18425;
squeal_samples[8183]=15303;
squeal_samples[8184]=12378;
squeal_samples[8185]=9648;
squeal_samples[8186]=7265;
squeal_samples[8187]=8890;
squeal_samples[8188]=11987;
squeal_samples[8189]=14977;
squeal_samples[8190]=17816;
squeal_samples[8191]=20553;
squeal_samples[8192]=23151;
squeal_samples[8193]=25654;
squeal_samples[8194]=28026;
squeal_samples[8195]=30310;
squeal_samples[8196]=32489;
squeal_samples[8197]=34576;
squeal_samples[8198]=36560;
squeal_samples[8199]=38459;
squeal_samples[8200]=40281;
squeal_samples[8201]=42012;
squeal_samples[8202]=43674;
squeal_samples[8203]=45255;
squeal_samples[8204]=46766;
squeal_samples[8205]=48212;
squeal_samples[8206]=49591;
squeal_samples[8207]=50913;
squeal_samples[8208]=51967;
squeal_samples[8209]=48482;
squeal_samples[8210]=43422;
squeal_samples[8211]=38698;
squeal_samples[8212]=34261;
squeal_samples[8213]=30124;
squeal_samples[8214]=26245;
squeal_samples[8215]=22623;
squeal_samples[8216]=19226;
squeal_samples[8217]=16049;
squeal_samples[8218]=13079;
squeal_samples[8219]=10301;
squeal_samples[8220]=7702;
squeal_samples[8221]=8078;
squeal_samples[8222]=11214;
squeal_samples[8223]=14225;
squeal_samples[8224]=17108;
squeal_samples[8225]=19862;
squeal_samples[8226]=22501;
squeal_samples[8227]=25025;
squeal_samples[8228]=27436;
squeal_samples[8229]=29735;
squeal_samples[8230]=31942;
squeal_samples[8231]=34043;
squeal_samples[8232]=36062;
squeal_samples[8233]=37980;
squeal_samples[8234]=39821;
squeal_samples[8235]=41574;
squeal_samples[8236]=43250;
squeal_samples[8237]=44853;
squeal_samples[8238]=46384;
squeal_samples[8239]=47845;
squeal_samples[8240]=49242;
squeal_samples[8241]=50574;
squeal_samples[8242]=51849;
squeal_samples[8243]=49785;
squeal_samples[8244]=44642;
squeal_samples[8245]=39836;
squeal_samples[8246]=35331;
squeal_samples[8247]=31120;
squeal_samples[8248]=27177;
squeal_samples[8249]=23496;
squeal_samples[8250]=20038;
squeal_samples[8251]=16807;
squeal_samples[8252]=13790;
squeal_samples[8253]=10960;
squeal_samples[8254]=8328;
squeal_samples[8255]=7438;
squeal_samples[8256]=10430;
squeal_samples[8257]=13473;
squeal_samples[8258]=16384;
squeal_samples[8259]=19177;
squeal_samples[8260]=21839;
squeal_samples[8261]=24397;
squeal_samples[8262]=26827;
squeal_samples[8263]=29163;
squeal_samples[8264]=31381;
squeal_samples[8265]=33520;
squeal_samples[8266]=35551;
squeal_samples[8267]=37496;
squeal_samples[8268]=39359;
squeal_samples[8269]=41129;
squeal_samples[8270]=42829;
squeal_samples[8271]=44441;
squeal_samples[8272]=45992;
squeal_samples[8273]=47473;
squeal_samples[8274]=48887;
squeal_samples[8275]=50234;
squeal_samples[8276]=51526;
squeal_samples[8277]=50903;
squeal_samples[8278]=45884;
squeal_samples[8279]=40998;
squeal_samples[8280]=36413;
squeal_samples[8281]=32135;
squeal_samples[8282]=28119;
squeal_samples[8283]=24380;
squeal_samples[8284]=20866;
squeal_samples[8285]=17583;
squeal_samples[8286]=14515;
squeal_samples[8287]=11638;
squeal_samples[8288]=8957;
squeal_samples[8289]=7147;
squeal_samples[8290]=9639;
squeal_samples[8291]=12711;
squeal_samples[8292]=15655;
squeal_samples[8293]=18473;
squeal_samples[8294]=21172;
squeal_samples[8295]=23750;
squeal_samples[8296]=26220;
squeal_samples[8297]=28572;
squeal_samples[8298]=30828;
squeal_samples[8299]=32979;
squeal_samples[8300]=35039;
squeal_samples[8301]=37006;
squeal_samples[8302]=38882;
squeal_samples[8303]=40680;
squeal_samples[8304]=42395;
squeal_samples[8305]=44032;
squeal_samples[8306]=45601;
squeal_samples[8307]=47092;
squeal_samples[8308]=48530;
squeal_samples[8309]=49886;
squeal_samples[8310]=51198;
squeal_samples[8311]=51975;
squeal_samples[8312]=47937;
squeal_samples[8313]=42912;
squeal_samples[8314]=38212;
squeal_samples[8315]=33812;
squeal_samples[8316]=29691;
squeal_samples[8317]=25844;
squeal_samples[8318]=22241;
squeal_samples[8319]=18868;
squeal_samples[8320]=15711;
squeal_samples[8321]=12763;
squeal_samples[8322]=10001;
squeal_samples[8323]=7468;
squeal_samples[8324]=8500;
squeal_samples[8325]=11622;
squeal_samples[8326]=14614;
squeal_samples[8327]=17478;
squeal_samples[8328]=20214;
squeal_samples[8329]=22835;
squeal_samples[8330]=25347;
squeal_samples[8331]=27730;
squeal_samples[8332]=30026;
squeal_samples[8333]=32215;
squeal_samples[8334]=34305;
squeal_samples[8335]=36309;
squeal_samples[8336]=38218;
squeal_samples[8337]=40043;
squeal_samples[8338]=41784;
squeal_samples[8339]=43451;
squeal_samples[8340]=45041;
squeal_samples[8341]=46563;
squeal_samples[8342]=48013;
squeal_samples[8343]=49397;
squeal_samples[8344]=50725;
squeal_samples[8345]=51995;
squeal_samples[8346]=49920;
squeal_samples[8347]=44767;
squeal_samples[8348]=39943;
squeal_samples[8349]=35433;
squeal_samples[8350]=31210;
squeal_samples[8351]=27266;
squeal_samples[8352]=23568;
squeal_samples[8353]=20110;
squeal_samples[8354]=16870;
squeal_samples[8355]=13849;
squeal_samples[8356]=11014;
squeal_samples[8357]=8371;
squeal_samples[8358]=7473;
squeal_samples[8359]=10469;
squeal_samples[8360]=13503;
squeal_samples[8361]=16417;
squeal_samples[8362]=19202;
squeal_samples[8363]=21862;
squeal_samples[8364]=24415;
squeal_samples[8365]=26851;
squeal_samples[8366]=29175;
squeal_samples[8367]=31399;
squeal_samples[8368]=33529;
squeal_samples[8369]=35560;
squeal_samples[8370]=37510;
squeal_samples[8371]=39357;
squeal_samples[8372]=41135;
squeal_samples[8373]=42822;
squeal_samples[8374]=44444;
squeal_samples[8375]=45990;
squeal_samples[8376]=47466;
squeal_samples[8377]=48881;
squeal_samples[8378]=50226;
squeal_samples[8379]=51516;
squeal_samples[8380]=51454;
squeal_samples[8381]=46651;
squeal_samples[8382]=41707;
squeal_samples[8383]=37076;
squeal_samples[8384]=32751;
squeal_samples[8385]=28699;
squeal_samples[8386]=24910;
squeal_samples[8387]=21370;
squeal_samples[8388]=18046;
squeal_samples[8389]=14949;
squeal_samples[8390]=12041;
squeal_samples[8391]=9328;
squeal_samples[8392]=7187;
squeal_samples[8393]=9279;
squeal_samples[8394]=12367;
squeal_samples[8395]=15329;
squeal_samples[8396]=18155;
squeal_samples[8397]=20869;
squeal_samples[8398]=23456;
squeal_samples[8399]=25938;
squeal_samples[8400]=28299;
squeal_samples[8401]=30567;
squeal_samples[8402]=32727;
squeal_samples[8403]=34796;
squeal_samples[8404]=36776;
squeal_samples[8405]=38661;
squeal_samples[8406]=40465;
squeal_samples[8407]=42190;
squeal_samples[8408]=43829;
squeal_samples[8409]=45410;
squeal_samples[8410]=46908;
squeal_samples[8411]=48348;
squeal_samples[8412]=49713;
squeal_samples[8413]=51027;
squeal_samples[8414]=52073;
squeal_samples[8415]=48577;
squeal_samples[8416]=43510;
squeal_samples[8417]=38764;
squeal_samples[8418]=34327;
squeal_samples[8419]=30175;
squeal_samples[8420]=26293;
squeal_samples[8421]=22661;
squeal_samples[8422]=19248;
squeal_samples[8423]=16074;
squeal_samples[8424]=13090;
squeal_samples[8425]=10312;
squeal_samples[8426]=7705;
squeal_samples[8427]=8077;
squeal_samples[8428]=11212;
squeal_samples[8429]=14219;
squeal_samples[8430]=17096;
squeal_samples[8431]=19853;
squeal_samples[8432]=22491;
squeal_samples[8433]=25005;
squeal_samples[8434]=27419;
squeal_samples[8435]=29713;
squeal_samples[8436]=31916;
squeal_samples[8437]=34024;
squeal_samples[8438]=36029;
squeal_samples[8439]=37954;
squeal_samples[8440]=39785;
squeal_samples[8441]=41540;
squeal_samples[8442]=43212;
squeal_samples[8443]=44812;
squeal_samples[8444]=46340;
squeal_samples[8445]=47799;
squeal_samples[8446]=49197;
squeal_samples[8447]=50528;
squeal_samples[8448]=51805;
squeal_samples[8449]=50499;
squeal_samples[8450]=45360;
squeal_samples[8451]=40495;
squeal_samples[8452]=35945;
squeal_samples[8453]=31686;
squeal_samples[8454]=27706;
squeal_samples[8455]=23980;
squeal_samples[8456]=20493;
squeal_samples[8457]=17231;
squeal_samples[8458]=14177;
squeal_samples[8459]=11320;
squeal_samples[8460]=8650;
squeal_samples[8461]=7259;
squeal_samples[8462]=10040;
squeal_samples[8463]=13098;
squeal_samples[8464]=16019;
squeal_samples[8465]=18820;
squeal_samples[8466]=21500;
squeal_samples[8467]=24064;
squeal_samples[8468]=26516;
squeal_samples[8469]=28852;
squeal_samples[8470]=31092;
squeal_samples[8471]=33225;
squeal_samples[8472]=35278;
squeal_samples[8473]=37225;
squeal_samples[8474]=39097;
squeal_samples[8475]=40875;
squeal_samples[8476]=42579;
squeal_samples[8477]=44210;
squeal_samples[8478]=45759;
squeal_samples[8479]=47251;
squeal_samples[8480]=48666;
squeal_samples[8481]=50022;
squeal_samples[8482]=51321;
squeal_samples[8483]=51727;
squeal_samples[8484]=47253;
squeal_samples[8485]=42272;
squeal_samples[8486]=37602;
squeal_samples[8487]=33240;
squeal_samples[8488]=29151;
squeal_samples[8489]=25337;
squeal_samples[8490]=21757;
squeal_samples[8491]=18412;
squeal_samples[8492]=15284;
squeal_samples[8493]=12355;
squeal_samples[8494]=9617;
squeal_samples[8495]=7233;
squeal_samples[8496]=8850;
squeal_samples[8497]=11955;
squeal_samples[8498]=14922;
squeal_samples[8499]=17775;
squeal_samples[8500]=20493;
squeal_samples[8501]=23107;
squeal_samples[8502]=25592;
squeal_samples[8503]=27973;
squeal_samples[8504]=30252;
squeal_samples[8505]=32429;
squeal_samples[8506]=34507;
squeal_samples[8507]=36493;
squeal_samples[8508]=38393;
squeal_samples[8509]=40205;
squeal_samples[8510]=41939;
squeal_samples[8511]=43590;
squeal_samples[8512]=45182;
squeal_samples[8513]=46683;
squeal_samples[8514]=48133;
squeal_samples[8515]=49502;
squeal_samples[8516]=50828;
squeal_samples[8517]=52032;
squeal_samples[8518]=49198;
squeal_samples[8519]=44083;
squeal_samples[8520]=39303;
squeal_samples[8521]=34825;
squeal_samples[8522]=30641;
squeal_samples[8523]=26729;
squeal_samples[8524]=23058;
squeal_samples[8525]=19633;
squeal_samples[8526]=16421;
squeal_samples[8527]=13418;
squeal_samples[8528]=10610;
squeal_samples[8529]=7988;
squeal_samples[8530]=7684;
squeal_samples[8531]=10788;
squeal_samples[8532]=13815;
squeal_samples[8533]=16704;
squeal_samples[8534]=19476;
squeal_samples[8535]=22122;
squeal_samples[8536]=24661;
squeal_samples[8537]=27084;
squeal_samples[8538]=29393;
squeal_samples[8539]=31606;
squeal_samples[8540]=33725;
squeal_samples[8541]=35746;
squeal_samples[8542]=37678;
squeal_samples[8543]=39515;
squeal_samples[8544]=41288;
squeal_samples[8545]=42963;
squeal_samples[8546]=44582;
squeal_samples[8547]=46114;
squeal_samples[8548]=47582;
squeal_samples[8549]=48985;
squeal_samples[8550]=50324;
squeal_samples[8551]=51610;
squeal_samples[8552]=50976;
squeal_samples[8553]=45952;
squeal_samples[8554]=41050;
squeal_samples[8555]=36458;
squeal_samples[8556]=32170;
squeal_samples[8557]=28150;
squeal_samples[8558]=24391;
squeal_samples[8559]=20882;
squeal_samples[8560]=17584;
squeal_samples[8561]=14513;
squeal_samples[8562]=11624;
squeal_samples[8563]=8941;
squeal_samples[8564]=7125;
squeal_samples[8565]=9613;
squeal_samples[8566]=12684;
squeal_samples[8567]=15620;
squeal_samples[8568]=18442;
squeal_samples[8569]=21131;
squeal_samples[8570]=23717;
squeal_samples[8571]=26173;
squeal_samples[8572]=28530;
squeal_samples[8573]=30772;
squeal_samples[8574]=32930;
squeal_samples[8575]=34988;
squeal_samples[8576]=36948;
squeal_samples[8577]=38831;
squeal_samples[8578]=40616;
squeal_samples[8579]=42338;
squeal_samples[8580]=43967;
squeal_samples[8581]=45535;
squeal_samples[8582]=47022;
squeal_samples[8583]=48457;
squeal_samples[8584]=49818;
squeal_samples[8585]=51119;
squeal_samples[8586]=51902;
squeal_samples[8587]=47860;
squeal_samples[8588]=42835;
squeal_samples[8589]=38131;
squeal_samples[8590]=33729;
squeal_samples[8591]=29612;
squeal_samples[8592]=25761;
squeal_samples[8593]=22156;
squeal_samples[8594]=18778;
squeal_samples[8595]=15627;
squeal_samples[8596]=12674;
squeal_samples[8597]=9915;
squeal_samples[8598]=7375;
squeal_samples[8599]=8413;
squeal_samples[8600]=11536;
squeal_samples[8601]=14521;
squeal_samples[8602]=17385;
squeal_samples[8603]=20122;
squeal_samples[8604]=22744;
squeal_samples[8605]=25251;
squeal_samples[8606]=27642;
squeal_samples[8607]=29929;
squeal_samples[8608]=32121;
squeal_samples[8609]=34211;
squeal_samples[8610]=36212;
squeal_samples[8611]=38118;
squeal_samples[8612]=39947;
squeal_samples[8613]=41685;
squeal_samples[8614]=43355;
squeal_samples[8615]=44942;
squeal_samples[8616]=46464;
squeal_samples[8617]=47915;
squeal_samples[8618]=49300;
squeal_samples[8619]=50626;
squeal_samples[8620]=51898;
squeal_samples[8621]=50579;
squeal_samples[8622]=45434;
squeal_samples[8623]=40558;
squeal_samples[8624]=36007;
squeal_samples[8625]=31734;
squeal_samples[8626]=27745;
squeal_samples[8627]=24012;
squeal_samples[8628]=20524;
squeal_samples[8629]=17249;
squeal_samples[8630]=14197;
squeal_samples[8631]=11329;
squeal_samples[8632]=8658;
squeal_samples[8633]=7257;
squeal_samples[8634]=10039;
squeal_samples[8635]=13089;
squeal_samples[8636]=16017;
squeal_samples[8637]=18808;
squeal_samples[8638]=21490;
squeal_samples[8639]=24048;
squeal_samples[8640]=26501;
squeal_samples[8641]=28829;
squeal_samples[8642]=31072;
squeal_samples[8643]=33205;
squeal_samples[8644]=35254;
squeal_samples[8645]=37202;
squeal_samples[8646]=39066;
squeal_samples[8647]=40852;
squeal_samples[8648]=42551;
squeal_samples[8649]=44177;
squeal_samples[8650]=45729;
squeal_samples[8651]=47212;
squeal_samples[8652]=48629;
squeal_samples[8653]=49986;
squeal_samples[8654]=51274;
squeal_samples[8655]=51694;
squeal_samples[8656]=47207;
squeal_samples[8657]=42230;
squeal_samples[8658]=37560;
squeal_samples[8659]=33195;
squeal_samples[8660]=29105;
squeal_samples[8661]=25288;
squeal_samples[8662]=21708;
squeal_samples[8663]=18364;
squeal_samples[8664]=15229;
squeal_samples[8665]=12303;
squeal_samples[8666]=9567;
squeal_samples[8667]=7181;
squeal_samples[8668]=8795;
squeal_samples[8669]=11900;
squeal_samples[8670]=14872;
squeal_samples[8671]=17716;
squeal_samples[8672]=20444;
squeal_samples[8673]=23049;
squeal_samples[8674]=25541;
squeal_samples[8675]=27914;
squeal_samples[8676]=30191;
squeal_samples[8677]=32370;
squeal_samples[8678]=34449;
squeal_samples[8679]=36431;
squeal_samples[8680]=38338;
squeal_samples[8681]=40142;
squeal_samples[8682]=41880;
squeal_samples[8683]=43533;
squeal_samples[8684]=45114;
squeal_samples[8685]=46626;
squeal_samples[8686]=48072;
squeal_samples[8687]=49443;
squeal_samples[8688]=50768;
squeal_samples[8689]=52025;
squeal_samples[8690]=49946;
squeal_samples[8691]=44776;
squeal_samples[8692]=39951;
squeal_samples[8693]=35429;
squeal_samples[8694]=31199;
squeal_samples[8695]=27245;
squeal_samples[8696]=23544;
squeal_samples[8697]=20075;
squeal_samples[8698]=16838;
squeal_samples[8699]=13797;
squeal_samples[8700]=10962;
squeal_samples[8701]=8311;
squeal_samples[8702]=7417;
squeal_samples[8703]=10402;
squeal_samples[8704]=13442;
squeal_samples[8705]=16345;
squeal_samples[8706]=19127;
squeal_samples[8707]=21794;
squeal_samples[8708]=24338;
squeal_samples[8709]=26771;
squeal_samples[8710]=29095;
squeal_samples[8711]=31318;
squeal_samples[8712]=33443;
squeal_samples[8713]=35476;
squeal_samples[8714]=37414;
squeal_samples[8715]=39271;
squeal_samples[8716]=41040;
squeal_samples[8717]=42732;
squeal_samples[8718]=44352;
squeal_samples[8719]=45893;
squeal_samples[8720]=47369;
squeal_samples[8721]=48780;
squeal_samples[8722]=50123;
squeal_samples[8723]=51411;
squeal_samples[8724]=51816;
squeal_samples[8725]=47324;
squeal_samples[8726]=42333;
squeal_samples[8727]=37655;
squeal_samples[8728]=33281;
squeal_samples[8729]=29189;
squeal_samples[8730]=25363;
squeal_samples[8731]=21782;
squeal_samples[8732]=18423;
squeal_samples[8733]=15292;
squeal_samples[8734]=12356;
squeal_samples[8735]=9612;
squeal_samples[8736]=7226;
squeal_samples[8737]=8835;
squeal_samples[8738]=11932;
squeal_samples[8739]=14907;
squeal_samples[8740]=17743;
squeal_samples[8741]=20474;
squeal_samples[8742]=23070;
squeal_samples[8743]=25565;
squeal_samples[8744]=27935;
squeal_samples[8745]=30212;
squeal_samples[8746]=32384;
squeal_samples[8747]=34467;
squeal_samples[8748]=36445;
squeal_samples[8749]=38346;
squeal_samples[8750]=40159;
squeal_samples[8751]=41889;
squeal_samples[8752]=43540;
squeal_samples[8753]=45120;
squeal_samples[8754]=46630;
squeal_samples[8755]=48073;
squeal_samples[8756]=49451;
squeal_samples[8757]=50764;
squeal_samples[8758]=52024;
squeal_samples[8759]=49938;
squeal_samples[8760]=44775;
squeal_samples[8761]=39945;
squeal_samples[8762]=35426;
squeal_samples[8763]=31188;
squeal_samples[8764]=27236;
squeal_samples[8765]=23534;
squeal_samples[8766]=20060;
squeal_samples[8767]=16823;
squeal_samples[8768]=13786;
squeal_samples[8769]=10950;
squeal_samples[8770]=8293;
squeal_samples[8771]=7404;
squeal_samples[8772]=10385;
squeal_samples[8773]=13428;
squeal_samples[8774]=16330;
squeal_samples[8775]=19112;
squeal_samples[8776]=21773;
squeal_samples[8777]=24318;
squeal_samples[8778]=26756;
squeal_samples[8779]=29074;
squeal_samples[8780]=31299;
squeal_samples[8781]=33426;
squeal_samples[8782]=35457;
squeal_samples[8783]=37393;
squeal_samples[8784]=39250;
squeal_samples[8785]=41020;
squeal_samples[8786]=42712;
squeal_samples[8787]=44331;
squeal_samples[8788]=45872;
squeal_samples[8789]=47350;
squeal_samples[8790]=48757;
squeal_samples[8791]=50105;
squeal_samples[8792]=51389;
squeal_samples[8793]=51790;
squeal_samples[8794]=47304;
squeal_samples[8795]=42312;
squeal_samples[8796]=37634;
squeal_samples[8797]=33263;
squeal_samples[8798]=29165;
squeal_samples[8799]=25340;
squeal_samples[8800]=21753;
squeal_samples[8801]=18406;
squeal_samples[8802]=15263;
squeal_samples[8803]=12332;
squeal_samples[8804]=9586;
squeal_samples[8805]=7199;
squeal_samples[8806]=8810;
squeal_samples[8807]=11905;
squeal_samples[8808]=14882;
squeal_samples[8809]=17722;
squeal_samples[8810]=20449;
squeal_samples[8811]=23043;
squeal_samples[8812]=25541;
squeal_samples[8813]=27907;
squeal_samples[8814]=30186;
squeal_samples[8815]=32360;
squeal_samples[8816]=34439;
squeal_samples[8817]=36428;
squeal_samples[8818]=38316;
squeal_samples[8819]=40135;
squeal_samples[8820]=41863;
squeal_samples[8821]=43515;
squeal_samples[8822]=45093;
squeal_samples[8823]=46604;
squeal_samples[8824]=48047;
squeal_samples[8825]=49425;
squeal_samples[8826]=50739;
squeal_samples[8827]=51997;
squeal_samples[8828]=49914;
squeal_samples[8829]=44752;
squeal_samples[8830]=39921;
squeal_samples[8831]=35398;
squeal_samples[8832]=31170;
squeal_samples[8833]=27210;
squeal_samples[8834]=23505;
squeal_samples[8835]=20039;
squeal_samples[8836]=16792;
squeal_samples[8837]=13765;
squeal_samples[8838]=10920;
squeal_samples[8839]=8270;
squeal_samples[8840]=7374;
squeal_samples[8841]=10366;
squeal_samples[8842]=13395;
squeal_samples[8843]=16308;
squeal_samples[8844]=19085;
squeal_samples[8845]=21747;
squeal_samples[8846]=24293;
squeal_samples[8847]=26730;
squeal_samples[8848]=29047;
squeal_samples[8849]=31274;
squeal_samples[8850]=33399;
squeal_samples[8851]=35432;
squeal_samples[8852]=37367;
squeal_samples[8853]=39224;
squeal_samples[8854]=40993;
squeal_samples[8855]=42688;
squeal_samples[8856]=44303;
squeal_samples[8857]=45848;
squeal_samples[8858]=47323;
squeal_samples[8859]=48730;
squeal_samples[8860]=50081;
squeal_samples[8861]=51363;
squeal_samples[8862]=51763;
squeal_samples[8863]=47281;
squeal_samples[8864]=42282;
squeal_samples[8865]=37612;
squeal_samples[8866]=33233;
squeal_samples[8867]=29144;
squeal_samples[8868]=25311;
squeal_samples[8869]=21729;
squeal_samples[8870]=18378;
squeal_samples[8871]=15239;
squeal_samples[8872]=12304;
squeal_samples[8873]=9563;
squeal_samples[8874]=7170;
squeal_samples[8875]=8787;
squeal_samples[8876]=11877;
squeal_samples[8877]=14857;
squeal_samples[8878]=17696;
squeal_samples[8879]=20422;
squeal_samples[8880]=23019;
squeal_samples[8881]=25513;
squeal_samples[8882]=27883;
squeal_samples[8883]=30160;
squeal_samples[8884]=32332;
squeal_samples[8885]=34416;
squeal_samples[8886]=36398;
squeal_samples[8887]=38296;
squeal_samples[8888]=40104;
squeal_samples[8889]=41840;
squeal_samples[8890]=43487;
squeal_samples[8891]=45069;
squeal_samples[8892]=46577;
squeal_samples[8893]=48023;
squeal_samples[8894]=49396;
squeal_samples[8895]=50716;
squeal_samples[8896]=51970;
squeal_samples[8897]=49887;
squeal_samples[8898]=44728;
squeal_samples[8899]=39893;
squeal_samples[8900]=35374;
squeal_samples[8901]=31144;
squeal_samples[8902]=27182;
squeal_samples[8903]=23483;
squeal_samples[8904]=20007;
squeal_samples[8905]=16771;
squeal_samples[8906]=13737;
squeal_samples[8907]=10901;
squeal_samples[8908]=8243;
squeal_samples[8909]=7350;
squeal_samples[8910]=10335;
squeal_samples[8911]=13374;
squeal_samples[8912]=16280;
squeal_samples[8913]=19060;
squeal_samples[8914]=21720;
squeal_samples[8915]=24269;
squeal_samples[8916]=26700;
squeal_samples[8917]=29026;
squeal_samples[8918]=31244;
squeal_samples[8919]=33377;
squeal_samples[8920]=35403;
squeal_samples[8921]=37343;
squeal_samples[8922]=39197;
squeal_samples[8923]=40968;
squeal_samples[8924]=42661;
squeal_samples[8925]=44278;
squeal_samples[8926]=45822;
squeal_samples[8927]=47296;
squeal_samples[8928]=48707;
squeal_samples[8929]=50051;
squeal_samples[8930]=51339;
squeal_samples[8931]=51737;
squeal_samples[8932]=47255;
squeal_samples[8933]=42257;
squeal_samples[8934]=37584;
squeal_samples[8935]=33209;
squeal_samples[8936]=29115;
squeal_samples[8937]=25289;
squeal_samples[8938]=21700;
squeal_samples[8939]=18354;
squeal_samples[8940]=15210;
squeal_samples[8941]=12282;
squeal_samples[8942]=9533;
squeal_samples[8943]=7149;
squeal_samples[8944]=8755;
squeal_samples[8945]=11857;
squeal_samples[8946]=14826;
squeal_samples[8947]=17674;
squeal_samples[8948]=20393;
squeal_samples[8949]=22995;
squeal_samples[8950]=25486;
squeal_samples[8951]=27858;
squeal_samples[8952]=30132;
squeal_samples[8953]=32309;
squeal_samples[8954]=34386;
squeal_samples[8955]=36377;
squeal_samples[8956]=38263;
squeal_samples[8957]=40086;
squeal_samples[8958]=41806;
squeal_samples[8959]=43467;
squeal_samples[8960]=45039;
squeal_samples[8961]=46553;
squeal_samples[8962]=47995;
squeal_samples[8963]=49372;
squeal_samples[8964]=50685;
squeal_samples[8965]=51948;
squeal_samples[8966]=50624;
squeal_samples[8967]=45464;
squeal_samples[8968]=40584;
squeal_samples[8969]=36014;
squeal_samples[8970]=31743;
squeal_samples[8971]=27738;
squeal_samples[8972]=24003;
squeal_samples[8973]=20501;
squeal_samples[8974]=17219;
squeal_samples[8975]=14157;
squeal_samples[8976]=11294;
squeal_samples[8977]=8612;
squeal_samples[8978]=7213;
squeal_samples[8979]=9979;
squeal_samples[8980]=13036;
squeal_samples[8981]=15953;
squeal_samples[8982]=18746;
squeal_samples[8983]=21425;
squeal_samples[8984]=23978;
squeal_samples[8985]=26429;
squeal_samples[8986]=28757;
squeal_samples[8987]=30993;
squeal_samples[8988]=33126;
squeal_samples[8989]=35167;
squeal_samples[8990]=37120;
squeal_samples[8991]=38982;
squeal_samples[8992]=40762;
squeal_samples[8993]=42462;
squeal_samples[8994]=44084;
squeal_samples[8995]=45637;
squeal_samples[8996]=47120;
squeal_samples[8997]=48531;
squeal_samples[8998]=49887;
squeal_samples[8999]=51180;
squeal_samples[9000]=51952;
squeal_samples[9001]=47894;
squeal_samples[9002]=42860;
squeal_samples[9003]=38140;
squeal_samples[9004]=33735;
squeal_samples[9005]=29604;
squeal_samples[9006]=25744;
squeal_samples[9007]=22129;
squeal_samples[9008]=18741;
squeal_samples[9009]=15586;
squeal_samples[9010]=12621;
squeal_samples[9011]=9856;
squeal_samples[9012]=7315;
squeal_samples[9013]=8340;
squeal_samples[9014]=11464;
squeal_samples[9015]=14446;
squeal_samples[9016]=17305;
squeal_samples[9017]=20043;
squeal_samples[9018]=22659;
squeal_samples[9019]=25160;
squeal_samples[9020]=27552;
squeal_samples[9021]=29832;
squeal_samples[9022]=32025;
squeal_samples[9023]=34111;
squeal_samples[9024]=36108;
squeal_samples[9025]=38015;
squeal_samples[9026]=39836;
squeal_samples[9027]=41580;
squeal_samples[9028]=43242;
squeal_samples[9029]=44830;
squeal_samples[9030]=46346;
squeal_samples[9031]=47798;
squeal_samples[9032]=49178;
squeal_samples[9033]=50508;
squeal_samples[9034]=51768;
squeal_samples[9035]=51125;
squeal_samples[9036]=46071;
squeal_samples[9037]=41150;
squeal_samples[9038]=36549;
squeal_samples[9039]=32238;
squeal_samples[9040]=28200;
squeal_samples[9041]=24434;
squeal_samples[9042]=20898;
squeal_samples[9043]=17595;
squeal_samples[9044]=14506;
squeal_samples[9045]=11616;
squeal_samples[9046]=8912;
squeal_samples[9047]=7094;
squeal_samples[9048]=9569;
squeal_samples[9049]=12639;
squeal_samples[9050]=15568;
squeal_samples[9051]=18386;
squeal_samples[9052]=21069;
squeal_samples[9053]=23646;
squeal_samples[9054]=26103;
squeal_samples[9055]=28449;
squeal_samples[9056]=30696;
squeal_samples[9057]=32838;
squeal_samples[9058]=34898;
squeal_samples[9059]=36853;
squeal_samples[9060]=38732;
squeal_samples[9061]=40515;
squeal_samples[9062]=42232;
squeal_samples[9063]=43859;
squeal_samples[9064]=45424;
squeal_samples[9065]=46907;
squeal_samples[9066]=48340;
squeal_samples[9067]=49692;
squeal_samples[9068]=51000;
squeal_samples[9069]=52187;
squeal_samples[9070]=49328;
squeal_samples[9071]=44196;
squeal_samples[9072]=39391;
squeal_samples[9073]=34903;
squeal_samples[9074]=30691;
squeal_samples[9075]=26767;
squeal_samples[9076]=23078;
squeal_samples[9077]=19636;
squeal_samples[9078]=16410;
squeal_samples[9079]=13395;
squeal_samples[9080]=10580;
squeal_samples[9081]=7944;
squeal_samples[9082]=7627;
squeal_samples[9083]=10734;
squeal_samples[9084]=13748;
squeal_samples[9085]=16632;
squeal_samples[9086]=19397;
squeal_samples[9087]=22041;
squeal_samples[9088]=24571;
squeal_samples[9089]=26992;
squeal_samples[9090]=29293;
squeal_samples[9091]=31502;
squeal_samples[9092]=33613;
squeal_samples[9093]=35633;
squeal_samples[9094]=37558;
squeal_samples[9095]=39401;
squeal_samples[9096]=41155;
squeal_samples[9097]=42841;
squeal_samples[9098]=44447;
squeal_samples[9099]=45977;
squeal_samples[9100]=47445;
squeal_samples[9101]=48841;
squeal_samples[9102]=50178;
squeal_samples[9103]=51457;
squeal_samples[9104]=51851;
squeal_samples[9105]=47351;
squeal_samples[9106]=42347;
squeal_samples[9107]=37663;
squeal_samples[9108]=33282;
squeal_samples[9109]=29173;
squeal_samples[9110]=25342;
squeal_samples[9111]=21752;
squeal_samples[9112]=18389;
squeal_samples[9113]=15246;
squeal_samples[9114]=12307;
squeal_samples[9115]=9555;
squeal_samples[9116]=7166;
squeal_samples[9117]=8764;
squeal_samples[9118]=11870;
squeal_samples[9119]=14830;
squeal_samples[9120]=17675;
squeal_samples[9121]=20393;
squeal_samples[9122]=22994;
squeal_samples[9123]=25481;
squeal_samples[9124]=27853;
squeal_samples[9125]=30121;
squeal_samples[9126]=32292;
squeal_samples[9127]=34372;
squeal_samples[9128]=36352;
squeal_samples[9129]=38246;
squeal_samples[9130]=40058;
squeal_samples[9131]=41786;
squeal_samples[9132]=43440;
squeal_samples[9133]=45015;
squeal_samples[9134]=46525;
squeal_samples[9135]=47961;
squeal_samples[9136]=49342;
squeal_samples[9137]=50652;
squeal_samples[9138]=51915;
squeal_samples[9139]=50587;
squeal_samples[9140]=45426;
squeal_samples[9141]=40540;
squeal_samples[9142]=35972;
squeal_samples[9143]=31699;
squeal_samples[9144]=27694;
squeal_samples[9145]=23956;
squeal_samples[9146]=20451;
squeal_samples[9147]=17171;
squeal_samples[9148]=14109;
squeal_samples[9149]=11237;
squeal_samples[9150]=8561;
squeal_samples[9151]=7155;
squeal_samples[9152]=9930;
squeal_samples[9153]=12978;
squeal_samples[9154]=15901;
squeal_samples[9155]=18691;
squeal_samples[9156]=21370;
squeal_samples[9157]=23925;
squeal_samples[9158]=26370;
squeal_samples[9159]=28701;
squeal_samples[9160]=30942;
squeal_samples[9161]=33068;
squeal_samples[9162]=35116;
squeal_samples[9163]=37058;
squeal_samples[9164]=38925;
squeal_samples[9165]=40700;
squeal_samples[9166]=42404;
squeal_samples[9167]=44022;
squeal_samples[9168]=45580;
squeal_samples[9169]=47058;
squeal_samples[9170]=48474;
squeal_samples[9171]=49824;
squeal_samples[9172]=51122;
squeal_samples[9173]=52145;
squeal_samples[9174]=48631;
squeal_samples[9175]=43541;
squeal_samples[9176]=38779;
squeal_samples[9177]=34325;
squeal_samples[9178]=30153;
squeal_samples[9179]=26255;
squeal_samples[9180]=22599;
squeal_samples[9181]=19186;
squeal_samples[9182]=15982;
squeal_samples[9183]=13002;
squeal_samples[9184]=10194;
squeal_samples[9185]=7594;
squeal_samples[9186]=7944;
squeal_samples[9187]=11082;
squeal_samples[9188]=14078;
squeal_samples[9189]=16947;
squeal_samples[9190]=19700;
squeal_samples[9191]=22328;
squeal_samples[9192]=24840;
squeal_samples[9193]=27243;
squeal_samples[9194]=29534;
squeal_samples[9195]=31737;
squeal_samples[9196]=33833;
squeal_samples[9197]=35840;
squeal_samples[9198]=37756;
squeal_samples[9199]=39590;
squeal_samples[9200]=41335;
squeal_samples[9201]=43007;
squeal_samples[9202]=44604;
squeal_samples[9203]=46129;
squeal_samples[9204]=47584;
squeal_samples[9205]=48977;
squeal_samples[9206]=50306;
squeal_samples[9207]=51577;
squeal_samples[9208]=51497;
squeal_samples[9209]=46672;
squeal_samples[9210]=41704;
squeal_samples[9211]=37059;
squeal_samples[9212]=32716;
squeal_samples[9213]=28640;
squeal_samples[9214]=24842;
squeal_samples[9215]=21279;
squeal_samples[9216]=17948;
squeal_samples[9217]=14832;
squeal_samples[9218]=11914;
squeal_samples[9219]=9187;
squeal_samples[9220]=7036;
squeal_samples[9221]=9128;
squeal_samples[9222]=12201;
squeal_samples[9223]=15158;
squeal_samples[9224]=17982;
squeal_samples[9225]=20687;
squeal_samples[9226]=23269;
squeal_samples[9227]=25747;
squeal_samples[9228]=28101;
squeal_samples[9229]=30359;
squeal_samples[9230]=32520;
squeal_samples[9231]=34582;
squeal_samples[9232]=36557;
squeal_samples[9233]=38441;
squeal_samples[9234]=40237;
squeal_samples[9235]=41957;
squeal_samples[9236]=43603;
squeal_samples[9237]=45172;
squeal_samples[9238]=46669;
squeal_samples[9239]=48099;
squeal_samples[9240]=49469;
squeal_samples[9241]=50772;
squeal_samples[9242]=52029;
squeal_samples[9243]=49927;
squeal_samples[9244]=44758;
squeal_samples[9245]=39914;
squeal_samples[9246]=35386;
squeal_samples[9247]=31142;
squeal_samples[9248]=27174;
squeal_samples[9249]=23464;
squeal_samples[9250]=19990;
squeal_samples[9251]=16741;
squeal_samples[9252]=13700;
squeal_samples[9253]=10857;
squeal_samples[9254]=8201;
squeal_samples[9255]=7295;
squeal_samples[9256]=10283;
squeal_samples[9257]=13313;
squeal_samples[9258]=16216;
squeal_samples[9259]=18993;
squeal_samples[9260]=21660;
squeal_samples[9261]=24192;
squeal_samples[9262]=26631;
squeal_samples[9263]=28946;
squeal_samples[9264]=31170;
squeal_samples[9265]=33296;
squeal_samples[9266]=35321;
squeal_samples[9267]=37263;
squeal_samples[9268]=39108;
squeal_samples[9269]=40886;
squeal_samples[9270]=42563;
squeal_samples[9271]=44192;
squeal_samples[9272]=45725;
squeal_samples[9273]=47202;
squeal_samples[9274]=48607;
squeal_samples[9275]=49949;
squeal_samples[9276]=51241;
squeal_samples[9277]=51998;
squeal_samples[9278]=47938;
squeal_samples[9279]=42891;
squeal_samples[9280]=38167;
squeal_samples[9281]=33751;
squeal_samples[9282]=29606;
squeal_samples[9283]=25747;
squeal_samples[9284]=22117;
squeal_samples[9285]=18737;
squeal_samples[9286]=15561;
squeal_samples[9287]=12606;
squeal_samples[9288]=9823;
squeal_samples[9289]=7283;
squeal_samples[9290]=8303;
squeal_samples[9291]=11421;
squeal_samples[9292]=14407;
squeal_samples[9293]=17257;
squeal_samples[9294]=19995;
squeal_samples[9295]=22608;
squeal_samples[9296]=25111;
squeal_samples[9297]=27497;
squeal_samples[9298]=29778;
squeal_samples[9299]=31962;
squeal_samples[9300]=34052;
squeal_samples[9301]=36040;
squeal_samples[9302]=37957;
squeal_samples[9303]=39768;
squeal_samples[9304]=41512;
squeal_samples[9305]=43166;
squeal_samples[9306]=44761;
squeal_samples[9307]=46274;
squeal_samples[9308]=47725;
squeal_samples[9309]=49105;
squeal_samples[9310]=50426;
squeal_samples[9311]=51694;
squeal_samples[9312]=51606;
squeal_samples[9313]=46766;
squeal_samples[9314]=41797;
squeal_samples[9315]=37139;
squeal_samples[9316]=32786;
squeal_samples[9317]=28708;
squeal_samples[9318]=24910;
squeal_samples[9319]=21325;
squeal_samples[9320]=18004;
squeal_samples[9321]=14868;
squeal_samples[9322]=11955;
squeal_samples[9323]=9216;
squeal_samples[9324]=7064;
squeal_samples[9325]=9146;
squeal_samples[9326]=12229;
squeal_samples[9327]=15172;
squeal_samples[9328]=17998;
squeal_samples[9329]=20701;
squeal_samples[9330]=23280;
squeal_samples[9331]=25756;
squeal_samples[9332]=28111;
squeal_samples[9333]=30368;
squeal_samples[9334]=32526;
squeal_samples[9335]=34584;
squeal_samples[9336]=36558;
squeal_samples[9337]=38438;
squeal_samples[9338]=40238;
squeal_samples[9339]=41949;
squeal_samples[9340]=43597;
squeal_samples[9341]=45159;
squeal_samples[9342]=46657;
squeal_samples[9343]=48089;
squeal_samples[9344]=49454;
squeal_samples[9345]=50762;
squeal_samples[9346]=52007;
squeal_samples[9347]=50682;
squeal_samples[9348]=45501;
squeal_samples[9349]=40612;
squeal_samples[9350]=36027;
squeal_samples[9351]=31747;
squeal_samples[9352]=27737;
squeal_samples[9353]=23989;
squeal_samples[9354]=20478;
squeal_samples[9355]=17195;
squeal_samples[9356]=14123;
squeal_samples[9357]=11248;
squeal_samples[9358]=8563;
squeal_samples[9359]=7153;
squeal_samples[9360]=9929;
squeal_samples[9361]=12968;
squeal_samples[9362]=15891;
squeal_samples[9363]=18677;
squeal_samples[9364]=21351;
squeal_samples[9365]=23909;
squeal_samples[9366]=26348;
squeal_samples[9367]=28682;
squeal_samples[9368]=30908;
squeal_samples[9369]=33042;
squeal_samples[9370]=35079;
squeal_samples[9371]=37026;
squeal_samples[9372]=38888;
squeal_samples[9373]=40663;
squeal_samples[9374]=42359;
squeal_samples[9375]=43987;
squeal_samples[9376]=45531;
squeal_samples[9377]=47014;
squeal_samples[9378]=48428;
squeal_samples[9379]=49778;
squeal_samples[9380]=51071;
squeal_samples[9381]=52251;
squeal_samples[9382]=49382;
squeal_samples[9383]=44244;
squeal_samples[9384]=39425;
squeal_samples[9385]=34929;
squeal_samples[9386]=30707;
squeal_samples[9387]=26771;
squeal_samples[9388]=23079;
squeal_samples[9389]=19630;
squeal_samples[9390]=16393;
squeal_samples[9391]=13379;
squeal_samples[9392]=10547;
squeal_samples[9393]=7911;
squeal_samples[9394]=7585;
squeal_samples[9395]=10687;
squeal_samples[9396]=13702;
squeal_samples[9397]=16586;
squeal_samples[9398]=19345;
squeal_samples[9399]=21990;
squeal_samples[9400]=24513;
squeal_samples[9401]=26929;
squeal_samples[9402]=29236;
squeal_samples[9403]=31440;
squeal_samples[9404]=33550;
squeal_samples[9405]=35565;
squeal_samples[9406]=37491;
squeal_samples[9407]=39324;
squeal_samples[9408]=41086;
squeal_samples[9409]=42759;
squeal_samples[9410]=44368;
squeal_samples[9411]=45900;
squeal_samples[9412]=47359;
squeal_samples[9413]=48762;
squeal_samples[9414]=50093;
squeal_samples[9415]=51372;
squeal_samples[9416]=52125;
squeal_samples[9417]=48057;
squeal_samples[9418]=42991;
squeal_samples[9419]=38268;
squeal_samples[9420]=33828;
squeal_samples[9421]=29691;
squeal_samples[9422]=25808;
squeal_samples[9423]=22185;
squeal_samples[9424]=18787;
squeal_samples[9425]=15614;
squeal_samples[9426]=12638;
squeal_samples[9427]=9861;
squeal_samples[9428]=7304;
squeal_samples[9429]=8334;
squeal_samples[9430]=11435;
squeal_samples[9431]=14427;
squeal_samples[9432]=17271;
squeal_samples[9433]=20006;
squeal_samples[9434]=22618;
squeal_samples[9435]=25112;
squeal_samples[9436]=27499;
squeal_samples[9437]=29781;
squeal_samples[9438]=31964;
squeal_samples[9439]=34048;
squeal_samples[9440]=36040;
squeal_samples[9441]=37945;
squeal_samples[9442]=39762;
squeal_samples[9443]=41500;
squeal_samples[9444]=43161;
squeal_samples[9445]=44745;
squeal_samples[9446]=46257;
squeal_samples[9447]=47703;
squeal_samples[9448]=49087;
squeal_samples[9449]=50406;
squeal_samples[9450]=51670;
squeal_samples[9451]=51581;
squeal_samples[9452]=46741;
squeal_samples[9453]=41773;
squeal_samples[9454]=37112;
squeal_samples[9455]=32758;
squeal_samples[9456]=28678;
squeal_samples[9457]=24872;
squeal_samples[9458]=21299;
squeal_samples[9459]=17963;
squeal_samples[9460]=14832;
squeal_samples[9461]=11915;
squeal_samples[9462]=9184;
squeal_samples[9463]=7019;
squeal_samples[9464]=9110;
squeal_samples[9465]=12183;
squeal_samples[9466]=15136;
squeal_samples[9467]=17952;
squeal_samples[9468]=20659;
squeal_samples[9469]=23235;
squeal_samples[9470]=25714;
squeal_samples[9471]=28059;
squeal_samples[9472]=30329;
squeal_samples[9473]=32477;
squeal_samples[9474]=34545;
squeal_samples[9475]=36507;
squeal_samples[9476]=38394;
squeal_samples[9477]=40190;
squeal_samples[9478]=41909;
squeal_samples[9479]=43550;
squeal_samples[9480]=45113;
squeal_samples[9481]=46611;
squeal_samples[9482]=48042;
squeal_samples[9483]=49408;
squeal_samples[9484]=50715;
squeal_samples[9485]=51962;
squeal_samples[9486]=50633;
squeal_samples[9487]=45458;
squeal_samples[9488]=40563;
squeal_samples[9489]=35983;
squeal_samples[9490]=31699;
squeal_samples[9491]=27691;
squeal_samples[9492]=23943;
squeal_samples[9493]=20431;
squeal_samples[9494]=17145;
squeal_samples[9495]=14075;
squeal_samples[9496]=11202;
squeal_samples[9497]=8512;
squeal_samples[9498]=7099;
squeal_samples[9499]=9880;
squeal_samples[9500]=12920;
squeal_samples[9501]=15839;
squeal_samples[9502]=18627;
squeal_samples[9503]=21297;
squeal_samples[9504]=23858;
squeal_samples[9505]=26298;
squeal_samples[9506]=28626;
squeal_samples[9507]=30861;
squeal_samples[9508]=32988;
squeal_samples[9509]=35033;
squeal_samples[9510]=36975;
squeal_samples[9511]=38833;
squeal_samples[9512]=40621;
squeal_samples[9513]=42305;
squeal_samples[9514]=43937;
squeal_samples[9515]=45482;
squeal_samples[9516]=46964;
squeal_samples[9517]=48376;
squeal_samples[9518]=49726;
squeal_samples[9519]=51020;
squeal_samples[9520]=52198;
squeal_samples[9521]=49333;
squeal_samples[9522]=44188;
squeal_samples[9523]=39379;
squeal_samples[9524]=34871;
squeal_samples[9525]=30662;
squeal_samples[9526]=26720;
squeal_samples[9527]=23030;
squeal_samples[9528]=19576;
squeal_samples[9529]=16343;
squeal_samples[9530]=13327;
squeal_samples[9531]=10495;
squeal_samples[9532]=7859;
squeal_samples[9533]=7535;
squeal_samples[9534]=10638;
squeal_samples[9535]=13652;
squeal_samples[9536]=16534;
squeal_samples[9537]=19293;
squeal_samples[9538]=21938;
squeal_samples[9539]=24463;
squeal_samples[9540]=26874;
squeal_samples[9541]=29189;
squeal_samples[9542]=31384;
squeal_samples[9543]=33501;
squeal_samples[9544]=35512;
squeal_samples[9545]=37439;
squeal_samples[9546]=39274;
squeal_samples[9547]=41032;
squeal_samples[9548]=42709;
squeal_samples[9549]=44316;
squeal_samples[9550]=45848;
squeal_samples[9551]=47308;
squeal_samples[9552]=48709;
squeal_samples[9553]=50043;
squeal_samples[9554]=51317;
squeal_samples[9555]=52078;
squeal_samples[9556]=48000;
squeal_samples[9557]=42946;
squeal_samples[9558]=38209;
squeal_samples[9559]=33783;
squeal_samples[9560]=29632;
squeal_samples[9561]=25764;
squeal_samples[9562]=22127;
squeal_samples[9563]=18740;
squeal_samples[9564]=15559;
squeal_samples[9565]=12588;
squeal_samples[9566]=9808;
squeal_samples[9567]=7255;
squeal_samples[9568]=8278;
squeal_samples[9569]=11388;
squeal_samples[9570]=14371;
squeal_samples[9571]=17222;
squeal_samples[9572]=19954;
squeal_samples[9573]=22565;
squeal_samples[9574]=25061;
squeal_samples[9575]=27448;
squeal_samples[9576]=29727;
squeal_samples[9577]=31916;
squeal_samples[9578]=33994;
squeal_samples[9579]=35988;
squeal_samples[9580]=37894;
squeal_samples[9581]=39710;
squeal_samples[9582]=41449;
squeal_samples[9583]=43110;
squeal_samples[9584]=44691;
squeal_samples[9585]=46207;
squeal_samples[9586]=47651;
squeal_samples[9587]=49035;
squeal_samples[9588]=50356;
squeal_samples[9589]=51615;
squeal_samples[9590]=51533;
squeal_samples[9591]=46686;
squeal_samples[9592]=41723;
squeal_samples[9593]=37061;
squeal_samples[9594]=32705;
squeal_samples[9595]=28627;
squeal_samples[9596]=24819;
squeal_samples[9597]=21249;
squeal_samples[9598]=17910;
squeal_samples[9599]=14781;
squeal_samples[9600]=11864;
squeal_samples[9601]=9130;
squeal_samples[9602]=6971;
squeal_samples[9603]=9054;
squeal_samples[9604]=12135;
squeal_samples[9605]=15081;
squeal_samples[9606]=17904;
squeal_samples[9607]=20603;
squeal_samples[9608]=23189;
squeal_samples[9609]=25654;
squeal_samples[9610]=28018;
squeal_samples[9611]=30266;
squeal_samples[9612]=32435;
squeal_samples[9613]=34486;
squeal_samples[9614]=36459;
squeal_samples[9615]=38342;
squeal_samples[9616]=40137;
squeal_samples[9617]=41858;
squeal_samples[9618]=43499;
squeal_samples[9619]=45060;
squeal_samples[9620]=46561;
squeal_samples[9621]=47987;
squeal_samples[9622]=49359;
squeal_samples[9623]=50662;
squeal_samples[9624]=51911;
squeal_samples[9625]=50582;
squeal_samples[9626]=45403;
squeal_samples[9627]=40514;
squeal_samples[9628]=35930;
squeal_samples[9629]=31647;
squeal_samples[9630]=27641;
squeal_samples[9631]=23890;
squeal_samples[9632]=20379;
squeal_samples[9633]=17094;
squeal_samples[9634]=14022;
squeal_samples[9635]=11153;
squeal_samples[9636]=8457;
squeal_samples[9637]=7051;
squeal_samples[9638]=9824;
squeal_samples[9639]=12872;
squeal_samples[9640]=15785;
squeal_samples[9641]=18576;
squeal_samples[9642]=21245;
squeal_samples[9643]=23807;
squeal_samples[9644]=26245;
squeal_samples[9645]=28575;
squeal_samples[9646]=30809;
squeal_samples[9647]=32935;
squeal_samples[9648]=34984;
squeal_samples[9649]=36919;
squeal_samples[9650]=38787;
squeal_samples[9651]=40561;
squeal_samples[9652]=42262;
squeal_samples[9653]=43877;
squeal_samples[9654]=45437;
squeal_samples[9655]=46908;
squeal_samples[9656]=48324;
squeal_samples[9657]=49675;
squeal_samples[9658]=50966;
squeal_samples[9659]=52201;
squeal_samples[9660]=50091;
squeal_samples[9661]=44891;
squeal_samples[9662]=40037;
squeal_samples[9663]=35483;
squeal_samples[9664]=31227;
squeal_samples[9665]=27247;
squeal_samples[9666]=23519;
squeal_samples[9667]=20035;
squeal_samples[9668]=16769;
squeal_samples[9669]=13718;
squeal_samples[9670]=10866;
squeal_samples[9671]=8195;
squeal_samples[9672]=7282;
squeal_samples[9673]=10262;
squeal_samples[9674]=13288;
squeal_samples[9675]=16184;
squeal_samples[9676]=18960;
squeal_samples[9677]=21612;
squeal_samples[9678]=24152;
squeal_samples[9679]=26573;
squeal_samples[9680]=28897;
squeal_samples[9681]=31105;
squeal_samples[9682]=33232;
squeal_samples[9683]=35252;
squeal_samples[9684]=37189;
squeal_samples[9685]=39035;
squeal_samples[9686]=40804;
squeal_samples[9687]=42485;
squeal_samples[9688]=44099;
squeal_samples[9689]=45635;
squeal_samples[9690]=47111;
squeal_samples[9691]=48511;
squeal_samples[9692]=49852;
squeal_samples[9693]=51139;
squeal_samples[9694]=52307;
squeal_samples[9695]=49430;
squeal_samples[9696]=44277;
squeal_samples[9697]=39457;
squeal_samples[9698]=34946;
squeal_samples[9699]=30717;
squeal_samples[9700]=26773;
squeal_samples[9701]=23072;
squeal_samples[9702]=19614;
squeal_samples[9703]=16377;
squeal_samples[9704]=13351;
squeal_samples[9705]=10516;
squeal_samples[9706]=7866;
squeal_samples[9707]=7548;
squeal_samples[9708]=10643;
squeal_samples[9709]=13659;
squeal_samples[9710]=16532;
squeal_samples[9711]=19296;
squeal_samples[9712]=21929;
squeal_samples[9713]=24460;
squeal_samples[9714]=26864;
squeal_samples[9715]=29169;
squeal_samples[9716]=31373;
squeal_samples[9717]=33475;
squeal_samples[9718]=35494;
squeal_samples[9719]=37415;
squeal_samples[9720]=39253;
squeal_samples[9721]=41010;
squeal_samples[9722]=42683;
squeal_samples[9723]=44283;
squeal_samples[9724]=45815;
squeal_samples[9725]=47275;
squeal_samples[9726]=48673;
squeal_samples[9727]=50007;
squeal_samples[9728]=51284;
squeal_samples[9729]=52294;
squeal_samples[9730]=48760;
squeal_samples[9731]=43650;
squeal_samples[9732]=38862;
squeal_samples[9733]=34391;
squeal_samples[9734]=30197;
squeal_samples[9735]=26290;
squeal_samples[9736]=22617;
squeal_samples[9737]=19190;
squeal_samples[9738]=15977;
squeal_samples[9739]=12976;
squeal_samples[9740]=10164;
squeal_samples[9741]=7540;
squeal_samples[9742]=7891;
squeal_samples[9743]=11013;
squeal_samples[9744]=14009;
squeal_samples[9745]=16872;
squeal_samples[9746]=19620;
squeal_samples[9747]=22237;
squeal_samples[9748]=24754;
squeal_samples[9749]=27148;
squeal_samples[9750]=29435;
squeal_samples[9751]=31633;
squeal_samples[9752]=33722;
squeal_samples[9753]=35730;
squeal_samples[9754]=37637;
squeal_samples[9755]=39467;
squeal_samples[9756]=41209;
squeal_samples[9757]=42876;
squeal_samples[9758]=44471;
squeal_samples[9759]=45992;
squeal_samples[9760]=47442;
squeal_samples[9761]=48832;
squeal_samples[9762]=50159;
squeal_samples[9763]=51428;
squeal_samples[9764]=52167;
squeal_samples[9765]=48091;
squeal_samples[9766]=43015;
squeal_samples[9767]=38275;
squeal_samples[9768]=33840;
squeal_samples[9769]=29680;
squeal_samples[9770]=25803;
squeal_samples[9771]=22160;
squeal_samples[9772]=18763;
squeal_samples[9773]=15580;
squeal_samples[9774]=12597;
squeal_samples[9775]=9817;
squeal_samples[9776]=7252;
squeal_samples[9777]=8277;
squeal_samples[9778]=11385;
squeal_samples[9779]=14365;
squeal_samples[9780]=17208;
squeal_samples[9781]=19942;
squeal_samples[9782]=22546;
squeal_samples[9783]=25044;
squeal_samples[9784]=27428;
squeal_samples[9785]=29705;
squeal_samples[9786]=31885;
squeal_samples[9787]=33965;
squeal_samples[9788]=35961;
squeal_samples[9789]=37857;
squeal_samples[9790]=39677;
squeal_samples[9791]=41408;
squeal_samples[9792]=43069;
squeal_samples[9793]=44647;
squeal_samples[9794]=46165;
squeal_samples[9795]=47608;
squeal_samples[9796]=48987;
squeal_samples[9797]=50311;
squeal_samples[9798]=51563;
squeal_samples[9799]=51948;
squeal_samples[9800]=47421;
squeal_samples[9801]=42397;
squeal_samples[9802]=37690;
squeal_samples[9803]=33294;
squeal_samples[9804]=29169;
squeal_samples[9805]=25322;
squeal_samples[9806]=21713;
squeal_samples[9807]=18338;
squeal_samples[9808]=15179;
squeal_samples[9809]=12228;
squeal_samples[9810]=9464;
squeal_samples[9811]=7061;
squeal_samples[9812]=8662;
squeal_samples[9813]=11746;
squeal_samples[9814]=14715;
squeal_samples[9815]=17550;
squeal_samples[9816]=20258;
squeal_samples[9817]=22855;
squeal_samples[9818]=25335;
squeal_samples[9819]=27701;
squeal_samples[9820]=29971;
squeal_samples[9821]=32137;
squeal_samples[9822]=34207;
squeal_samples[9823]=36187;
squeal_samples[9824]=38077;
squeal_samples[9825]=39882;
squeal_samples[9826]=41606;
squeal_samples[9827]=43257;
squeal_samples[9828]=44831;
squeal_samples[9829]=46334;
squeal_samples[9830]=47771;
squeal_samples[9831]=49141;
squeal_samples[9832]=50457;
squeal_samples[9833]=51709;
squeal_samples[9834]=51612;
squeal_samples[9835]=46763;
squeal_samples[9836]=41779;
squeal_samples[9837]=37115;
squeal_samples[9838]=32747;
squeal_samples[9839]=28662;
squeal_samples[9840]=24848;
squeal_samples[9841]=21265;
squeal_samples[9842]=17918;
squeal_samples[9843]=14787;
squeal_samples[9844]=11860;
squeal_samples[9845]=9121;
squeal_samples[9846]=6961;
squeal_samples[9847]=9039;
squeal_samples[9848]=12115;
squeal_samples[9849]=15060;
squeal_samples[9850]=17879;
squeal_samples[9851]=20577;
squeal_samples[9852]=23155;
squeal_samples[9853]=25627;
squeal_samples[9854]=27976;
squeal_samples[9855]=30235;
squeal_samples[9856]=32389;
squeal_samples[9857]=34445;
squeal_samples[9858]=36417;
squeal_samples[9859]=38292;
squeal_samples[9860]=40093;
squeal_samples[9861]=41802;
squeal_samples[9862]=43447;
squeal_samples[9863]=45007;
squeal_samples[9864]=46507;
squeal_samples[9865]=47935;
squeal_samples[9866]=49299;
squeal_samples[9867]=50604;
squeal_samples[9868]=51852;
squeal_samples[9869]=51178;
squeal_samples[9870]=46111;
squeal_samples[9871]=41160;
squeal_samples[9872]=36545;
squeal_samples[9873]=32205;
squeal_samples[9874]=28158;
squeal_samples[9875]=24370;
squeal_samples[9876]=20821;
squeal_samples[9877]=17498;
squeal_samples[9878]=14404;
squeal_samples[9879]=11491;
squeal_samples[9880]=8783;
squeal_samples[9881]=6948;
squeal_samples[9882]=9417;
squeal_samples[9883]=12477;
squeal_samples[9884]=15406;
squeal_samples[9885]=18206;
squeal_samples[9886]=20897;
squeal_samples[9887]=23458;
squeal_samples[9888]=25910;
squeal_samples[9889]=28253;
squeal_samples[9890]=30491;
squeal_samples[9891]=32638;
squeal_samples[9892]=34681;
squeal_samples[9893]=36643;
squeal_samples[9894]=38507;
squeal_samples[9895]=40297;
squeal_samples[9896]=41995;
squeal_samples[9897]=43635;
squeal_samples[9898]=45183;
squeal_samples[9899]=46675;
squeal_samples[9900]=48095;
squeal_samples[9901]=49449;
squeal_samples[9902]=50749;
squeal_samples[9903]=51990;
squeal_samples[9904]=50647;
squeal_samples[9905]=45457;
squeal_samples[9906]=40562;
squeal_samples[9907]=35965;
squeal_samples[9908]=31678;
squeal_samples[9909]=27649;
squeal_samples[9910]=23906;
squeal_samples[9911]=20381;
squeal_samples[9912]=17092;
squeal_samples[9913]=14014;
squeal_samples[9914]=11130;
squeal_samples[9915]=8439;
squeal_samples[9916]=7020;
squeal_samples[9917]=9798;
squeal_samples[9918]=12837;
squeal_samples[9919]=15753;
squeal_samples[9920]=18534;
squeal_samples[9921]=21210;
squeal_samples[9922]=23759;
squeal_samples[9923]=26197;
squeal_samples[9924]=28526;
squeal_samples[9925]=30757;
squeal_samples[9926]=32882;
squeal_samples[9927]=34922;
squeal_samples[9928]=36864;
squeal_samples[9929]=38726;
squeal_samples[9930]=40498;
squeal_samples[9931]=42195;
squeal_samples[9932]=43818;
squeal_samples[9933]=45359;
squeal_samples[9934]=46842;
squeal_samples[9935]=48249;
squeal_samples[9936]=49605;
squeal_samples[9937]=50894;
squeal_samples[9938]=52125;
squeal_samples[9939]=50013;
squeal_samples[9940]=44814;
squeal_samples[9941]=39955;
squeal_samples[9942]=35401;
squeal_samples[9943]=31146;
squeal_samples[9944]=27156;
squeal_samples[9945]=23434;
squeal_samples[9946]=19944;
squeal_samples[9947]=16685;
squeal_samples[9948]=13628;
squeal_samples[9949]=10774;
squeal_samples[9950]=8101;
squeal_samples[9951]=7189;
squeal_samples[9952]=10169;
squeal_samples[9953]=13194;
squeal_samples[9954]=16093;
squeal_samples[9955]=18863;
squeal_samples[9956]=21524;
squeal_samples[9957]=24053;
squeal_samples[9958]=26485;
squeal_samples[9959]=28793;
squeal_samples[9960]=31015;
squeal_samples[9961]=33132;
squeal_samples[9962]=35154;
squeal_samples[9963]=37090;
squeal_samples[9964]=38936;
squeal_samples[9965]=40703;
squeal_samples[9966]=42390;
squeal_samples[9967]=44002;
squeal_samples[9968]=45539;
squeal_samples[9969]=47011;
squeal_samples[9970]=48411;
squeal_samples[9971]=49754;
squeal_samples[9972]=51038;
squeal_samples[9973]=52263;
squeal_samples[9974]=50141;
squeal_samples[9975]=44933;
squeal_samples[9976]=40065;
squeal_samples[9977]=35508;
squeal_samples[9978]=31239;
squeal_samples[9979]=27248;
squeal_samples[9980]=23517;
squeal_samples[9981]=20021;
squeal_samples[9982]=16749;
squeal_samples[9983]=13695;
squeal_samples[9984]=10832;
squeal_samples[9985]=8157;
squeal_samples[9986]=7238;
squeal_samples[9987]=10218;
squeal_samples[9988]=13240;
squeal_samples[9989]=16138;
squeal_samples[9990]=18906;
squeal_samples[9991]=21558;
squeal_samples[9992]=24090;
squeal_samples[9993]=26521;
squeal_samples[9994]=28827;
squeal_samples[9995]=31048;
squeal_samples[9996]=33159;
squeal_samples[9997]=35182;
squeal_samples[9998]=37112;
squeal_samples[9999]=38964;
squeal_samples[10000]=40722;
squeal_samples[10001]=42408;
squeal_samples[10002]=44018;
squeal_samples[10003]=45551;
squeal_samples[10004]=47027;
squeal_samples[10005]=48425;
squeal_samples[10006]=49769;
squeal_samples[10007]=51046;
squeal_samples[10008]=52225;
squeal_samples[10009]=49339;
squeal_samples[10010]=44186;
squeal_samples[10011]=39364;
squeal_samples[10012]=34846;
squeal_samples[10013]=30626;
squeal_samples[10014]=26674;
squeal_samples[10015]=22973;
squeal_samples[10016]=19512;
squeal_samples[10017]=16277;
squeal_samples[10018]=13243;
squeal_samples[10019]=10417;
squeal_samples[10020]=7763;
squeal_samples[10021]=7442;
squeal_samples[10022]=10538;
squeal_samples[10023]=13550;
squeal_samples[10024]=16429;
squeal_samples[10025]=19186;
squeal_samples[10026]=21826;
squeal_samples[10027]=24349;
squeal_samples[10028]=26763;
squeal_samples[10029]=29058;
squeal_samples[10030]=31269;
squeal_samples[10031]=33367;
squeal_samples[10032]=35388;
squeal_samples[10033]=37303;
squeal_samples[10034]=39141;
squeal_samples[10035]=40898;
squeal_samples[10036]=42575;
squeal_samples[10037]=44179;
squeal_samples[10038]=45700;
squeal_samples[10039]=47166;
squeal_samples[10040]=48557;
squeal_samples[10041]=49897;
squeal_samples[10042]=51171;
squeal_samples[10043]=52333;
squeal_samples[10044]=49448;
squeal_samples[10045]=44286;
squeal_samples[10046]=39457;
squeal_samples[10047]=34936;
squeal_samples[10048]=30699;
squeal_samples[10049]=26752;
squeal_samples[10050]=23044;
squeal_samples[10051]=19576;
squeal_samples[10052]=16334;
squeal_samples[10053]=13302;
squeal_samples[10054]=10460;
squeal_samples[10055]=7813;
squeal_samples[10056]=7485;
squeal_samples[10057]=10582;
squeal_samples[10058]=13584;
squeal_samples[10059]=16464;
squeal_samples[10060]=19218;
squeal_samples[10061]=21854;
squeal_samples[10062]=24377;
squeal_samples[10063]=26783;
squeal_samples[10064]=29088;
squeal_samples[10065]=31289;
squeal_samples[10066]=33391;
squeal_samples[10067]=35404;
squeal_samples[10068]=37324;
squeal_samples[10069]=39160;
squeal_samples[10070]=40912;
squeal_samples[10071]=42590;
squeal_samples[10072]=44190;
squeal_samples[10073]=45718;
squeal_samples[10074]=47176;
squeal_samples[10075]=48573;
squeal_samples[10076]=49907;
squeal_samples[10077]=51174;
squeal_samples[10078]=52349;
squeal_samples[10079]=49450;
squeal_samples[10080]=44292;
squeal_samples[10081]=39461;
squeal_samples[10082]=34935;
squeal_samples[10083]=30707;
squeal_samples[10084]=26746;
squeal_samples[10085]=23043;
squeal_samples[10086]=19574;
squeal_samples[10087]=16330;
squeal_samples[10088]=13301;
squeal_samples[10089]=10457;
squeal_samples[10090]=7806;
squeal_samples[10091]=7477;
squeal_samples[10092]=10574;
squeal_samples[10093]=13575;
squeal_samples[10094]=16459;
squeal_samples[10095]=19212;
squeal_samples[10096]=21850;
squeal_samples[10097]=24372;
squeal_samples[10098]=26782;
squeal_samples[10099]=29079;
squeal_samples[10100]=31282;
squeal_samples[10101]=33383;
squeal_samples[10102]=35396;
squeal_samples[10103]=37317;
squeal_samples[10104]=39151;
squeal_samples[10105]=40906;
squeal_samples[10106]=42580;
squeal_samples[10107]=44180;
squeal_samples[10108]=45706;
squeal_samples[10109]=47171;
squeal_samples[10110]=48560;
squeal_samples[10111]=49897;
squeal_samples[10112]=51171;
squeal_samples[10113]=52335;
squeal_samples[10114]=49447;
squeal_samples[10115]=44282;
squeal_samples[10116]=39448;
squeal_samples[10117]=34928;
squeal_samples[10118]=30694;
squeal_samples[10119]=26737;
squeal_samples[10120]=23033;
squeal_samples[10121]=19561;
squeal_samples[10122]=16322;
squeal_samples[10123]=13284;
squeal_samples[10124]=10451;
squeal_samples[10125]=7799;
squeal_samples[10126]=7462;
squeal_samples[10127]=10562;
squeal_samples[10128]=13567;
squeal_samples[10129]=16451;
squeal_samples[10130]=19198;
squeal_samples[10131]=21839;
squeal_samples[10132]=24356;
squeal_samples[10133]=26772;
squeal_samples[10134]=29064;
squeal_samples[10135]=31269;
squeal_samples[10136]=33375;
squeal_samples[10137]=35383;
squeal_samples[10138]=37303;
squeal_samples[10139]=39140;
squeal_samples[10140]=40889;
squeal_samples[10141]=42571;
squeal_samples[10142]=44163;
squeal_samples[10143]=45696;
squeal_samples[10144]=47156;
squeal_samples[10145]=48553;
squeal_samples[10146]=49883;
squeal_samples[10147]=51157;
squeal_samples[10148]=52324;
squeal_samples[10149]=49432;
squeal_samples[10150]=44270;
squeal_samples[10151]=39434;
squeal_samples[10152]=34915;
squeal_samples[10153]=30679;
squeal_samples[10154]=26727;
squeal_samples[10155]=23015;
squeal_samples[10156]=19554;
squeal_samples[10157]=16303;
squeal_samples[10158]=13274;
squeal_samples[10159]=10437;
squeal_samples[10160]=7785;
squeal_samples[10161]=7450;
squeal_samples[10162]=10548;
squeal_samples[10163]=13554;
squeal_samples[10164]=16438;
squeal_samples[10165]=19185;
squeal_samples[10166]=21830;
squeal_samples[10167]=24343;
squeal_samples[10168]=26759;
squeal_samples[10169]=29051;
squeal_samples[10170]=31256;
squeal_samples[10171]=33362;
squeal_samples[10172]=35368;
squeal_samples[10173]=37292;
squeal_samples[10174]=39124;
squeal_samples[10175]=40879;
squeal_samples[10176]=42555;
squeal_samples[10177]=44151;
squeal_samples[10178]=45683;
squeal_samples[10179]=47141;
squeal_samples[10180]=48542;
squeal_samples[10181]=49867;
squeal_samples[10182]=51147;
squeal_samples[10183]=52308;
squeal_samples[10184]=49421;
squeal_samples[10185]=44255;
squeal_samples[10186]=39422;
squeal_samples[10187]=34901;
squeal_samples[10188]=30666;
squeal_samples[10189]=26714;
squeal_samples[10190]=23002;
squeal_samples[10191]=19540;
squeal_samples[10192]=16291;
squeal_samples[10193]=13259;
squeal_samples[10194]=10426;
squeal_samples[10195]=7769;
squeal_samples[10196]=7440;
squeal_samples[10197]=10531;
squeal_samples[10198]=13545;
squeal_samples[10199]=16420;
squeal_samples[10200]=19177;
squeal_samples[10201]=21813;
squeal_samples[10202]=24332;
squeal_samples[10203]=26745;
squeal_samples[10204]=29036;
squeal_samples[10205]=31246;
squeal_samples[10206]=33345;
squeal_samples[10207]=35359;
squeal_samples[10208]=37274;
squeal_samples[10209]=39116;
squeal_samples[10210]=40861;
squeal_samples[10211]=42545;
squeal_samples[10212]=44136;
squeal_samples[10213]=45668;
squeal_samples[10214]=47132;
squeal_samples[10215]=48524;
squeal_samples[10216]=49859;
squeal_samples[10217]=51128;
squeal_samples[10218]=52300;
squeal_samples[10219]=49402;
squeal_samples[10220]=44247;
squeal_samples[10221]=39404;
squeal_samples[10222]=34892;
squeal_samples[10223]=30650;
squeal_samples[10224]=26702;
squeal_samples[10225]=22988;
squeal_samples[10226]=19526;
squeal_samples[10227]=16279;
squeal_samples[10228]=13245;
squeal_samples[10229]=10413;
squeal_samples[10230]=7756;
squeal_samples[10231]=7425;
squeal_samples[10232]=10521;
squeal_samples[10233]=13528;
squeal_samples[10234]=16410;
squeal_samples[10235]=19160;
squeal_samples[10236]=21802;
squeal_samples[10237]=24318;
squeal_samples[10238]=26732;
squeal_samples[10239]=29023;
squeal_samples[10240]=31230;
squeal_samples[10241]=33335;
squeal_samples[10242]=35342;
squeal_samples[10243]=37266;
squeal_samples[10244]=39097;
squeal_samples[10245]=40851;
squeal_samples[10246]=42530;
squeal_samples[10247]=44123;
squeal_samples[10248]=45658;
squeal_samples[10249]=47115;
squeal_samples[10250]=48512;
squeal_samples[10251]=49845;
squeal_samples[10252]=51116;
squeal_samples[10253]=52285;
squeal_samples[10254]=49391;
squeal_samples[10255]=44231;
squeal_samples[10256]=39393;
squeal_samples[10257]=34877;
squeal_samples[10258]=30639;
squeal_samples[10259]=26684;
squeal_samples[10260]=22980;
squeal_samples[10261]=19509;
squeal_samples[10262]=16268;
squeal_samples[10263]=13231;
squeal_samples[10264]=10399;
squeal_samples[10265]=7743;
squeal_samples[10266]=7412;
squeal_samples[10267]=10508;
squeal_samples[10268]=13513;
squeal_samples[10269]=16399;
squeal_samples[10270]=19145;
squeal_samples[10271]=21789;
squeal_samples[10272]=24306;
squeal_samples[10273]=26716;
squeal_samples[10274]=29013;
squeal_samples[10275]=31215;
squeal_samples[10276]=33321;
squeal_samples[10277]=35331;
squeal_samples[10278]=37249;
squeal_samples[10279]=39088;
squeal_samples[10280]=40835;
squeal_samples[10281]=42517;
squeal_samples[10282]=44110;
squeal_samples[10283]=45644;
squeal_samples[10284]=47101;
squeal_samples[10285]=48502;
squeal_samples[10286]=49827;
squeal_samples[10287]=51107;
squeal_samples[10288]=52267;
squeal_samples[10289]=49382;
squeal_samples[10290]=44214;
squeal_samples[10291]=39384;
squeal_samples[10292]=34859;
squeal_samples[10293]=30628;
squeal_samples[10294]=26671;
squeal_samples[10295]=22964;
squeal_samples[10296]=19500;
squeal_samples[10297]=16250;
squeal_samples[10298]=13220;
squeal_samples[10299]=10385;
squeal_samples[10300]=7729;
squeal_samples[10301]=7401;
squeal_samples[10302]=10491;
squeal_samples[10303]=13503;
squeal_samples[10304]=16381;
squeal_samples[10305]=19136;
squeal_samples[10306]=21774;
squeal_samples[10307]=24292;
squeal_samples[10308]=26704;
squeal_samples[10309]=28996;
squeal_samples[10310]=31205;
squeal_samples[10311]=33306;
squeal_samples[10312]=35319;
squeal_samples[10313]=37234;
squeal_samples[10314]=39073;
squeal_samples[10315]=40825;
squeal_samples[10316]=42499;
squeal_samples[10317]=44103;
squeal_samples[10318]=45623;
squeal_samples[10319]=47093;
squeal_samples[10320]=48483;
squeal_samples[10321]=49818;
squeal_samples[10322]=51089;
squeal_samples[10323]=52306;
squeal_samples[10324]=50173;
squeal_samples[10325]=44961;
squeal_samples[10326]=40075;
squeal_samples[10327]=35516;
squeal_samples[10328]=31231;
squeal_samples[10329]=27239;
squeal_samples[10330]=23496;
squeal_samples[10331]=19997;
squeal_samples[10332]=16715;
squeal_samples[10333]=13652;
squeal_samples[10334]=10783;
squeal_samples[10335]=8104;
squeal_samples[10336]=7183;
squeal_samples[10337]=10158;
squeal_samples[10338]=13180;
squeal_samples[10339]=16070;
squeal_samples[10340]=18838;
squeal_samples[10341]=21484;
squeal_samples[10342]=24018;
squeal_samples[10343]=26440;
squeal_samples[10344]=28751;
squeal_samples[10345]=30963;
squeal_samples[10346]=33074;
squeal_samples[10347]=35100;
squeal_samples[10348]=37025;
squeal_samples[10349]=38871;
squeal_samples[10350]=40629;
squeal_samples[10351]=42318;
squeal_samples[10352]=43917;
squeal_samples[10353]=45462;
squeal_samples[10354]=46920;
squeal_samples[10355]=48328;
squeal_samples[10356]=49660;
squeal_samples[10357]=50946;
squeal_samples[10358]=52165;
squeal_samples[10359]=50811;
squeal_samples[10360]=45599;
squeal_samples[10361]=40682;
squeal_samples[10362]=36065;
squeal_samples[10363]=31757;
squeal_samples[10364]=27720;
squeal_samples[10365]=23953;
squeal_samples[10366]=20415;
squeal_samples[10367]=17117;
squeal_samples[10368]=14021;
squeal_samples[10369]=11131;
squeal_samples[10370]=8425;
squeal_samples[10371]=7003;
squeal_samples[10372]=9764;
squeal_samples[10373]=12800;
squeal_samples[10374]=15712;
squeal_samples[10375]=18490;
squeal_samples[10376]=21160;
squeal_samples[10377]=23695;
squeal_samples[10378]=26143;
squeal_samples[10379]=28459;
squeal_samples[10380]=30683;
squeal_samples[10381]=32809;
squeal_samples[10382]=34836;
squeal_samples[10383]=36785;
squeal_samples[10384]=38633;
squeal_samples[10385]=40412;
squeal_samples[10386]=42095;
squeal_samples[10387]=43722;
squeal_samples[10388]=45257;
squeal_samples[10389]=46737;
squeal_samples[10390]=48144;
squeal_samples[10391]=49489;
squeal_samples[10392]=50781;
squeal_samples[10393]=52009;
squeal_samples[10394]=51324;
squeal_samples[10395]=46229;
squeal_samples[10396]=41263;
squeal_samples[10397]=36619;
squeal_samples[10398]=32269;
squeal_samples[10399]=28201;
squeal_samples[10400]=24401;
squeal_samples[10401]=20836;
squeal_samples[10402]=17503;
squeal_samples[10403]=14387;
squeal_samples[10404]=11467;
squeal_samples[10405]=8746;
squeal_samples[10406]=6900;
squeal_samples[10407]=9365;
squeal_samples[10408]=12419;
squeal_samples[10409]=15342;
squeal_samples[10410]=18138;
squeal_samples[10411]=20817;
squeal_samples[10412]=23377;
squeal_samples[10413]=25827;
squeal_samples[10414]=28159;
squeal_samples[10415]=30397;
squeal_samples[10416]=32536;
squeal_samples[10417]=34580;
squeal_samples[10418]=36529;
squeal_samples[10419]=38396;
squeal_samples[10420]=40176;
squeal_samples[10421]=41881;
squeal_samples[10422]=43503;
squeal_samples[10423]=45056;
squeal_samples[10424]=46544;
squeal_samples[10425]=47961;
squeal_samples[10426]=49314;
squeal_samples[10427]=50609;
squeal_samples[10428]=51842;
squeal_samples[10429]=51731;
squeal_samples[10430]=46854;
squeal_samples[10431]=41856;
squeal_samples[10432]=37168;
squeal_samples[10433]=32788;
squeal_samples[10434]=28683;
squeal_samples[10435]=24846;
squeal_samples[10436]=21261;
squeal_samples[10437]=17895;
squeal_samples[10438]=14753;
squeal_samples[10439]=11813;
squeal_samples[10440]=9064;
squeal_samples[10441]=6885;
squeal_samples[10442]=8963;
squeal_samples[10443]=12028;
squeal_samples[10444]=14971;
squeal_samples[10445]=17783;
squeal_samples[10446]=20475;
squeal_samples[10447]=23052;
squeal_samples[10448]=25512;
squeal_samples[10449]=27861;
squeal_samples[10450]=30110;
squeal_samples[10451]=32262;
squeal_samples[10452]=34317;
squeal_samples[10453]=36277;
squeal_samples[10454]=38154;
squeal_samples[10455]=39946;
squeal_samples[10456]=41656;
squeal_samples[10457]=43292;
squeal_samples[10458]=44856;
squeal_samples[10459]=46342;
squeal_samples[10460]=47776;
squeal_samples[10461]=49132;
squeal_samples[10462]=50436;
squeal_samples[10463]=51680;
squeal_samples[10464]=52032;
squeal_samples[10465]=47498;
squeal_samples[10466]=42446;
squeal_samples[10467]=37729;
squeal_samples[10468]=33306;
squeal_samples[10469]=29166;
squeal_samples[10470]=25304;
squeal_samples[10471]=21676;
squeal_samples[10472]=18294;
squeal_samples[10473]=15117;
squeal_samples[10474]=12153;
squeal_samples[10475]=9382;
squeal_samples[10476]=6965;
squeal_samples[10477]=8556;
squeal_samples[10478]=11641;
squeal_samples[10479]=14599;
squeal_samples[10480]=17426;
squeal_samples[10481]=20133;
squeal_samples[10482]=22720;
squeal_samples[10483]=25198;
squeal_samples[10484]=27556;
squeal_samples[10485]=29824;
squeal_samples[10486]=31984;
squeal_samples[10487]=34052;
squeal_samples[10488]=36021;
squeal_samples[10489]=37916;
squeal_samples[10490]=39712;
squeal_samples[10491]=41438;
squeal_samples[10492]=43079;
squeal_samples[10493]=44649;
squeal_samples[10494]=46153;
squeal_samples[10495]=47585;
squeal_samples[10496]=48957;
squeal_samples[10497]=50260;
squeal_samples[10498]=51512;
squeal_samples[10499]=52238;
squeal_samples[10500]=48134;
squeal_samples[10501]=43048;
squeal_samples[10502]=38285;
squeal_samples[10503]=33829;
squeal_samples[10504]=29656;
squeal_samples[10505]=25758;
squeal_samples[10506]=22107;
squeal_samples[10507]=18689;
squeal_samples[10508]=15491;
squeal_samples[10509]=12505;
squeal_samples[10510]=9702;
squeal_samples[10511]=7135;
squeal_samples[10512]=8143;
squeal_samples[10513]=11246;
squeal_samples[10514]=14225;
squeal_samples[10515]=17061;
squeal_samples[10516]=19791;
squeal_samples[10517]=22390;
squeal_samples[10518]=24880;
squeal_samples[10519]=27257;
squeal_samples[10520]=29531;
squeal_samples[10521]=31706;
squeal_samples[10522]=33787;
squeal_samples[10523]=35771;
squeal_samples[10524]=37668;
squeal_samples[10525]=39477;
squeal_samples[10526]=41211;
squeal_samples[10527]=42865;
squeal_samples[10528]=44446;
squeal_samples[10529]=45954;
squeal_samples[10530]=47395;
squeal_samples[10531]=48771;
squeal_samples[10532]=50092;
squeal_samples[10533]=51343;
squeal_samples[10534]=52340;
squeal_samples[10535]=48784;
squeal_samples[10536]=43654;
squeal_samples[10537]=38851;
squeal_samples[10538]=34356;
squeal_samples[10539]=30147;
squeal_samples[10540]=26225;
squeal_samples[10541]=22532;
squeal_samples[10542]=19092;
squeal_samples[10543]=15863;
squeal_samples[10544]=12846;
squeal_samples[10545]=10032;
squeal_samples[10546]=7386;
squeal_samples[10547]=7736;
squeal_samples[10548]=10853;
squeal_samples[10549]=13844;
squeal_samples[10550]=16698;
squeal_samples[10551]=19444;
squeal_samples[10552]=22055;
squeal_samples[10553]=24566;
squeal_samples[10554]=26945;
squeal_samples[10555]=29245;
squeal_samples[10556]=31425;
squeal_samples[10557]=33518;
squeal_samples[10558]=35514;
squeal_samples[10559]=37419;
squeal_samples[10560]=39242;
squeal_samples[10561]=40987;
squeal_samples[10562]=42644;
squeal_samples[10563]=44237;
squeal_samples[10564]=45756;
squeal_samples[10565]=47205;
squeal_samples[10566]=48594;
squeal_samples[10567]=49910;
squeal_samples[10568]=51182;
squeal_samples[10569]=52332;
squeal_samples[10570]=49437;
squeal_samples[10571]=44256;
squeal_samples[10572]=39423;
squeal_samples[10573]=34886;
squeal_samples[10574]=30650;
squeal_samples[10575]=26677;
squeal_samples[10576]=22968;
squeal_samples[10577]=19496;
squeal_samples[10578]=16237;
squeal_samples[10579]=13207;
squeal_samples[10580]=10355;
squeal_samples[10581]=7699;
squeal_samples[10582]=7367;
squeal_samples[10583]=10458;
squeal_samples[10584]=13461;
squeal_samples[10585]=16338;
squeal_samples[10586]=19091;
squeal_samples[10587]=21726;
squeal_samples[10588]=24244;
squeal_samples[10589]=26647;
squeal_samples[10590]=28947;
squeal_samples[10591]=31140;
squeal_samples[10592]=33250;
squeal_samples[10593]=35256;
squeal_samples[10594]=37172;
squeal_samples[10595]=39006;
squeal_samples[10596]=40760;
squeal_samples[10597]=42432;
squeal_samples[10598]=44024;
squeal_samples[10599]=45557;
squeal_samples[10600]=47009;
squeal_samples[10601]=48407;
squeal_samples[10602]=49735;
squeal_samples[10603]=51007;
squeal_samples[10604]=52229;
squeal_samples[10605]=50095;
squeal_samples[10606]=44875;
squeal_samples[10607]=39993;
squeal_samples[10608]=35424;
squeal_samples[10609]=31143;
squeal_samples[10610]=27151;
squeal_samples[10611]=23401;
squeal_samples[10612]=19909;
squeal_samples[10613]=16617;
squeal_samples[10614]=13565;
squeal_samples[10615]=10687;
squeal_samples[10616]=8014;
squeal_samples[10617]=7084;
squeal_samples[10618]=10060;
squeal_samples[10619]=13084;
squeal_samples[10620]=15969;
squeal_samples[10621]=18744;
squeal_samples[10622]=21383;
squeal_samples[10623]=23922;
squeal_samples[10624]=26342;
squeal_samples[10625]=28647;
squeal_samples[10626]=30865;
squeal_samples[10627]=32972;
squeal_samples[10628]=34994;
squeal_samples[10629]=36925;
squeal_samples[10630]=38769;
squeal_samples[10631]=40530;
squeal_samples[10632]=42211;
squeal_samples[10633]=43816;
squeal_samples[10634]=45356;
squeal_samples[10635]=46819;
squeal_samples[10636]=48222;
squeal_samples[10637]=49559;
squeal_samples[10638]=50839;
squeal_samples[10639]=52064;
squeal_samples[10640]=51368;
squeal_samples[10641]=46262;
squeal_samples[10642]=41297;
squeal_samples[10643]=36638;
squeal_samples[10644]=32292;
squeal_samples[10645]=28207;
squeal_samples[10646]=24401;
squeal_samples[10647]=20831;
squeal_samples[10648]=17492;
squeal_samples[10649]=14375;
squeal_samples[10650]=11445;
squeal_samples[10651]=8718;
squeal_samples[10652]=6867;
squeal_samples[10653]=9337;
squeal_samples[10654]=12382;
squeal_samples[10655]=15301;
squeal_samples[10656]=18097;
squeal_samples[10657]=20775;
squeal_samples[10658]=23330;
squeal_samples[10659]=25782;
squeal_samples[10660]=28111;
squeal_samples[10661]=30348;
squeal_samples[10662]=32479;
squeal_samples[10663]=34525;
squeal_samples[10664]=36472;
squeal_samples[10665]=38337;
squeal_samples[10666]=40122;
squeal_samples[10667]=41814;
squeal_samples[10668]=43442;
squeal_samples[10669]=44992;
squeal_samples[10670]=46476;
squeal_samples[10671]=47893;
squeal_samples[10672]=49246;
squeal_samples[10673]=50534;
squeal_samples[10674]=51769;
squeal_samples[10675]=51661;
squeal_samples[10676]=46782;
squeal_samples[10677]=41780;
squeal_samples[10678]=37091;
squeal_samples[10679]=32707;
squeal_samples[10680]=28603;
squeal_samples[10681]=24769;
squeal_samples[10682]=21172;
squeal_samples[10683]=17814;
squeal_samples[10684]=14665;
squeal_samples[10685]=11730;
squeal_samples[10686]=8975;
squeal_samples[10687]=7114;
squeal_samples[10688]=9563;
squeal_samples[10689]=12604;
squeal_samples[10690]=15515;
squeal_samples[10691]=18299;
squeal_samples[10692]=20969;
squeal_samples[10693]=23512;
squeal_samples[10694]=25949;
squeal_samples[10695]=28282;
squeal_samples[10696]=30501;
squeal_samples[10697]=32635;
squeal_samples[10698]=34665;
squeal_samples[10699]=36610;
squeal_samples[10700]=38466;
squeal_samples[10701]=40242;
squeal_samples[10702]=41931;
squeal_samples[10703]=43554;
squeal_samples[10704]=45097;
squeal_samples[10705]=46577;
squeal_samples[10706]=47986;
squeal_samples[10707]=49337;
squeal_samples[10708]=50621;
squeal_samples[10709]=51858;
squeal_samples[10710]=51729;
squeal_samples[10711]=46859;
squeal_samples[10712]=41839;
squeal_samples[10713]=37155;
squeal_samples[10714]=32765;
squeal_samples[10715]=28653;
squeal_samples[10716]=24816;
squeal_samples[10717]=21218;
squeal_samples[10718]=17854;
squeal_samples[10719]=14703;
squeal_samples[10720]=11756;
squeal_samples[10721]=9011;
squeal_samples[10722]=6828;
squeal_samples[10723]=8904;
squeal_samples[10724]=11967;
squeal_samples[10725]=14905;
squeal_samples[10726]=17717;
squeal_samples[10727]=20403;
squeal_samples[10728]=22981;
squeal_samples[10729]=25442;
squeal_samples[10730]=27786;
squeal_samples[10731]=30037;
squeal_samples[10732]=32182;
squeal_samples[10733]=34236;
squeal_samples[10734]=36201;
squeal_samples[10735]=38071;
squeal_samples[10736]=39863;
squeal_samples[10737]=41574;
squeal_samples[10738]=43205;
squeal_samples[10739]=44771;
squeal_samples[10740]=46257;
squeal_samples[10741]=47687;
squeal_samples[10742]=49044;
squeal_samples[10743]=50343;
squeal_samples[10744]=51590;
squeal_samples[10745]=52304;
squeal_samples[10746]=48192;
squeal_samples[10747]=43093;
squeal_samples[10748]=38323;
squeal_samples[10749]=33861;
squeal_samples[10750]=29674;
squeal_samples[10751]=25777;
squeal_samples[10752]=22109;
squeal_samples[10753]=18689;
squeal_samples[10754]=15486;
squeal_samples[10755]=12488;
squeal_samples[10756]=9686;
squeal_samples[10757]=7112;
squeal_samples[10758]=8118;
squeal_samples[10759]=11218;
squeal_samples[10760]=14188;
squeal_samples[10761]=17032;
squeal_samples[10762]=19748;
squeal_samples[10763]=22354;
squeal_samples[10764]=24834;
squeal_samples[10765]=27212;
squeal_samples[10766]=29482;
squeal_samples[10767]=31656;
squeal_samples[10768]=33732;
squeal_samples[10769]=35715;
squeal_samples[10770]=37613;
squeal_samples[10771]=39421;
squeal_samples[10772]=41151;
squeal_samples[10773]=42804;
squeal_samples[10774]=44379;
squeal_samples[10775]=45894;
squeal_samples[10776]=47327;
squeal_samples[10777]=48707;
squeal_samples[10778]=50018;
squeal_samples[10779]=51276;
squeal_samples[10780]=52428;
squeal_samples[10781]=49513;
squeal_samples[10782]=44330;
squeal_samples[10783]=39477;
squeal_samples[10784]=34937;
squeal_samples[10785]=30690;
squeal_samples[10786]=26710;
squeal_samples[10787]=22994;
squeal_samples[10788]=19516;
squeal_samples[10789]=16253;
squeal_samples[10790]=13210;
squeal_samples[10791]=10360;
squeal_samples[10792]=7697;
squeal_samples[10793]=7360;
squeal_samples[10794]=10448;
squeal_samples[10795]=13447;
squeal_samples[10796]=16321;
squeal_samples[10797]=19069;
squeal_samples[10798]=21702;
squeal_samples[10799]=24215;
squeal_samples[10800]=26617;
squeal_samples[10801]=28913;
squeal_samples[10802]=31112;
squeal_samples[10803]=33207;
squeal_samples[10804]=35219;
squeal_samples[10805]=37131;
squeal_samples[10806]=38969;
squeal_samples[10807]=40714;
squeal_samples[10808]=42387;
squeal_samples[10809]=43983;
squeal_samples[10810]=45506;
squeal_samples[10811]=46965;
squeal_samples[10812]=48353;
squeal_samples[10813]=49685;
squeal_samples[10814]=50958;
squeal_samples[10815]=52173;
squeal_samples[10816]=50799;
squeal_samples[10817]=45581;
squeal_samples[10818]=40649;
squeal_samples[10819]=36030;
squeal_samples[10820]=31715;
squeal_samples[10821]=27667;
squeal_samples[10822]=23889;
squeal_samples[10823]=20346;
squeal_samples[10824]=17036;
squeal_samples[10825]=13937;
squeal_samples[10826]=11045;
squeal_samples[10827]=8329;
squeal_samples[10828]=6901;
squeal_samples[10829]=9662;
squeal_samples[10830]=12693;
squeal_samples[10831]=15605;
squeal_samples[10832]=18377;
squeal_samples[10833]=21047;
squeal_samples[10834]=23579;
squeal_samples[10835]=26017;
squeal_samples[10836]=28338;
squeal_samples[10837]=30557;
squeal_samples[10838]=32681;
squeal_samples[10839]=34708;
squeal_samples[10840]=36649;
squeal_samples[10841]=38501;
squeal_samples[10842]=40275;
squeal_samples[10843]=41957;
squeal_samples[10844]=43580;
squeal_samples[10845]=45118;
squeal_samples[10846]=46592;
squeal_samples[10847]=47998;
squeal_samples[10848]=49344;
squeal_samples[10849]=50629;
squeal_samples[10850]=51858;
squeal_samples[10851]=51738;
squeal_samples[10852]=46855;
squeal_samples[10853]=41841;
squeal_samples[10854]=37146;
squeal_samples[10855]=32754;
squeal_samples[10856]=28642;
squeal_samples[10857]=24798;
squeal_samples[10858]=21196;
squeal_samples[10859]=17831;
squeal_samples[10860]=14680;
squeal_samples[10861]=11735;
squeal_samples[10862]=8981;
squeal_samples[10863]=6797;
squeal_samples[10864]=8874;
squeal_samples[10865]=11934;
squeal_samples[10866]=14873;
squeal_samples[10867]=17681;
squeal_samples[10868]=20373;
squeal_samples[10869]=22946;
squeal_samples[10870]=25402;
squeal_samples[10871]=27751;
squeal_samples[10872]=29993;
squeal_samples[10873]=32148;
squeal_samples[10874]=34194;
squeal_samples[10875]=36163;
squeal_samples[10876]=38033;
squeal_samples[10877]=39824;
squeal_samples[10878]=41534;
squeal_samples[10879]=43168;
squeal_samples[10880]=44724;
squeal_samples[10881]=46216;
squeal_samples[10882]=47640;
squeal_samples[10883]=49000;
squeal_samples[10884]=50300;
squeal_samples[10885]=51538;
squeal_samples[10886]=52262;
squeal_samples[10887]=48146;
squeal_samples[10888]=43049;
squeal_samples[10889]=38274;
squeal_samples[10890]=33810;
squeal_samples[10891]=29627;
squeal_samples[10892]=25723;
squeal_samples[10893]=22064;
squeal_samples[10894]=18634;
squeal_samples[10895]=15436;
squeal_samples[10896]=12435;
squeal_samples[10897]=9638;
squeal_samples[10898]=7061;
squeal_samples[10899]=8069;
squeal_samples[10900]=11168;
squeal_samples[10901]=14133;
squeal_samples[10902]=16981;
squeal_samples[10903]=19695;
squeal_samples[10904]=22302;
squeal_samples[10905]=24787;
squeal_samples[10906]=27159;
squeal_samples[10907]=29435;
squeal_samples[10908]=31605;
squeal_samples[10909]=33677;
squeal_samples[10910]=35665;
squeal_samples[10911]=37557;
squeal_samples[10912]=39373;
squeal_samples[10913]=41095;
squeal_samples[10914]=42755;
squeal_samples[10915]=44322;
squeal_samples[10916]=45840;
squeal_samples[10917]=47272;
squeal_samples[10918]=48651;
squeal_samples[10919]=49963;
squeal_samples[10920]=51223;
squeal_samples[10921]=52369;
squeal_samples[10922]=49461;
squeal_samples[10923]=44278;
squeal_samples[10924]=39423;
squeal_samples[10925]=34883;
squeal_samples[10926]=30633;
squeal_samples[10927]=26661;
squeal_samples[10928]=22939;
squeal_samples[10929]=19460;
squeal_samples[10930]=16200;
squeal_samples[10931]=13153;
squeal_samples[10932]=10305;
squeal_samples[10933]=7644;
squeal_samples[10934]=7301;
squeal_samples[10935]=10396;
squeal_samples[10936]=13391;
squeal_samples[10937]=16266;
squeal_samples[10938]=19013;
squeal_samples[10939]=21647;
squeal_samples[10940]=24160;
squeal_samples[10941]=26562;
squeal_samples[10942]=28859;
squeal_samples[10943]=31054;
squeal_samples[10944]=33154;
squeal_samples[10945]=35162;
squeal_samples[10946]=37078;
squeal_samples[10947]=38913;
squeal_samples[10948]=40658;
squeal_samples[10949]=42332;
squeal_samples[10950]=43927;
squeal_samples[10951]=45452;
squeal_samples[10952]=46909;
squeal_samples[10953]=48298;
squeal_samples[10954]=49629;
squeal_samples[10955]=50903;
squeal_samples[10956]=52117;
squeal_samples[10957]=50744;
squeal_samples[10958]=45527;
squeal_samples[10959]=40592;
squeal_samples[10960]=35975;
squeal_samples[10961]=31660;
squeal_samples[10962]=27610;
squeal_samples[10963]=23835;
squeal_samples[10964]=20290;
squeal_samples[10965]=16980;
squeal_samples[10966]=13883;
squeal_samples[10967]=10987;
squeal_samples[10968]=8275;
squeal_samples[10969]=7331;
squeal_samples[10970]=10289;
squeal_samples[10971]=13289;
squeal_samples[10972]=16172;
squeal_samples[10973]=18922;
squeal_samples[10974]=21557;
squeal_samples[10975]=24076;
squeal_samples[10976]=26481;
squeal_samples[10977]=28782;
squeal_samples[10978]=30979;
squeal_samples[10979]=33082;
squeal_samples[10980]=35086;
squeal_samples[10981]=37012;
squeal_samples[10982]=38843;
squeal_samples[10983]=40596;
squeal_samples[10984]=42270;
squeal_samples[10985]=43863;
squeal_samples[10986]=45396;
squeal_samples[10987]=46850;
squeal_samples[10988]=48247;
squeal_samples[10989]=49577;
squeal_samples[10990]=50851;
squeal_samples[10991]=52064;
squeal_samples[10992]=51366;
squeal_samples[10993]=46257;
squeal_samples[10994]=41274;
squeal_samples[10995]=36614;
squeal_samples[10996]=32253;
squeal_samples[10997]=28167;
squeal_samples[10998]=24354;
squeal_samples[10999]=20774;
squeal_samples[11000]=17437;
squeal_samples[11001]=14300;
squeal_samples[11002]=11384;
squeal_samples[11003]=8640;
squeal_samples[11004]=6795;
squeal_samples[11005]=9247;
squeal_samples[11006]=12304;
squeal_samples[11007]=15212;
squeal_samples[11008]=18019;
squeal_samples[11009]=20681;
squeal_samples[11010]=23245;
squeal_samples[11011]=25683;
squeal_samples[11012]=28016;
squeal_samples[11013]=30249;
squeal_samples[11014]=32382;
squeal_samples[11015]=34425;
squeal_samples[11016]=36369;
squeal_samples[11017]=38236;
squeal_samples[11018]=40011;
squeal_samples[11019]=41713;
squeal_samples[11020]=43334;
squeal_samples[11021]=44883;
squeal_samples[11022]=46363;
squeal_samples[11023]=47778;
squeal_samples[11024]=49126;
squeal_samples[11025]=50426;
squeal_samples[11026]=51654;
squeal_samples[11027]=52373;
squeal_samples[11028]=48239;
squeal_samples[11029]=43138;
squeal_samples[11030]=38351;
squeal_samples[11031]=33881;
squeal_samples[11032]=29690;
squeal_samples[11033]=25778;
squeal_samples[11034]=22110;
squeal_samples[11035]=18678;
squeal_samples[11036]=15471;
squeal_samples[11037]=12462;
squeal_samples[11038]=9664;
squeal_samples[11039]=7074;
squeal_samples[11040]=8088;
squeal_samples[11041]=11175;
squeal_samples[11042]=14144;
squeal_samples[11043]=16985;
squeal_samples[11044]=19698;
squeal_samples[11045]=22302;
squeal_samples[11046]=24787;
squeal_samples[11047]=27152;
squeal_samples[11048]=29427;
squeal_samples[11049]=31594;
squeal_samples[11050]=33670;
squeal_samples[11051]=35654;
squeal_samples[11052]=37540;
squeal_samples[11053]=39354;
squeal_samples[11054]=41078;
squeal_samples[11055]=42731;
squeal_samples[11056]=44308;
squeal_samples[11057]=45813;
squeal_samples[11058]=47251;
squeal_samples[11059]=48628;
squeal_samples[11060]=49939;
squeal_samples[11061]=51194;
squeal_samples[11062]=52396;
squeal_samples[11063]=50239;
squeal_samples[11064]=45003;
squeal_samples[11065]=40098;
squeal_samples[11066]=35518;
squeal_samples[11067]=31219;
squeal_samples[11068]=27202;
squeal_samples[11069]=23449;
squeal_samples[11070]=19930;
squeal_samples[11071]=16639;
squeal_samples[11072]=13560;
squeal_samples[11073]=10679;
squeal_samples[11074]=7989;
squeal_samples[11075]=7059;
squeal_samples[11076]=10021;
squeal_samples[11077]=13039;
squeal_samples[11078]=15922;
squeal_samples[11079]=18686;
squeal_samples[11080]=21327;
squeal_samples[11081]=23854;
squeal_samples[11082]=26271;
squeal_samples[11083]=28573;
squeal_samples[11084]=30780;
squeal_samples[11085]=32893;
squeal_samples[11086]=34906;
squeal_samples[11087]=36832;
squeal_samples[11088]=38672;
squeal_samples[11089]=40431;
squeal_samples[11090]=42106;
squeal_samples[11091]=43717;
squeal_samples[11092]=45243;
squeal_samples[11093]=46707;
squeal_samples[11094]=48105;
squeal_samples[11095]=49441;
squeal_samples[11096]=50714;
squeal_samples[11097]=51938;
squeal_samples[11098]=51806;
squeal_samples[11099]=46916;
squeal_samples[11100]=41892;
squeal_samples[11101]=37184;
squeal_samples[11102]=32783;
squeal_samples[11103]=28664;
squeal_samples[11104]=24814;
squeal_samples[11105]=21210;
squeal_samples[11106]=17830;
squeal_samples[11107]=14676;
squeal_samples[11108]=11724;
squeal_samples[11109]=8967;
squeal_samples[11110]=6776;
squeal_samples[11111]=8847;
squeal_samples[11112]=11908;
squeal_samples[11113]=14846;
squeal_samples[11114]=17649;
squeal_samples[11115]=20338;
squeal_samples[11116]=22904;
squeal_samples[11117]=25365;
squeal_samples[11118]=27704;
squeal_samples[11119]=29953;
squeal_samples[11120]=32098;
squeal_samples[11121]=34148;
squeal_samples[11122]=36108;
squeal_samples[11123]=37980;
squeal_samples[11124]=39764;
squeal_samples[11125]=41477;
squeal_samples[11126]=43102;
squeal_samples[11127]=44662;
squeal_samples[11128]=46154;
squeal_samples[11129]=47577;
squeal_samples[11130]=48936;
squeal_samples[11131]=50234;
squeal_samples[11132]=51475;
squeal_samples[11133]=52451;
squeal_samples[11134]=48877;
squeal_samples[11135]=43721;
squeal_samples[11136]=38902;
squeal_samples[11137]=34384;
squeal_samples[11138]=30167;
squeal_samples[11139]=26217;
squeal_samples[11140]=22522;
squeal_samples[11141]=19058;
squeal_samples[11142]=15827;
squeal_samples[11143]=12790;
squeal_samples[11144]=9963;
squeal_samples[11145]=7315;
squeal_samples[11146]=7648;
squeal_samples[11147]=10765;
squeal_samples[11148]=13738;
squeal_samples[11149]=16601;
squeal_samples[11150]=19323;
squeal_samples[11151]=21946;
squeal_samples[11152]=24441;
squeal_samples[11153]=26822;
squeal_samples[11154]=29111;
squeal_samples[11155]=31290;
squeal_samples[11156]=33375;
squeal_samples[11157]=35367;
squeal_samples[11158]=37271;
squeal_samples[11159]=39089;
squeal_samples[11160]=40827;
squeal_samples[11161]=42487;
squeal_samples[11162]=44072;
squeal_samples[11163]=45587;
squeal_samples[11164]=47035;
squeal_samples[11165]=48418;
squeal_samples[11166]=49735;
squeal_samples[11167]=51000;
squeal_samples[11168]=52207;
squeal_samples[11169]=50829;
squeal_samples[11170]=45602;
squeal_samples[11171]=40655;
squeal_samples[11172]=36029;
squeal_samples[11173]=31700;
squeal_samples[11174]=27648;
squeal_samples[11175]=23865;
squeal_samples[11176]=20316;
squeal_samples[11177]=16997;
squeal_samples[11178]=13890;
squeal_samples[11179]=10987;
squeal_samples[11180]=8274;
squeal_samples[11181]=6835;
squeal_samples[11182]=9599;
squeal_samples[11183]=12622;
squeal_samples[11184]=15533;
squeal_samples[11185]=18299;
squeal_samples[11186]=20966;
squeal_samples[11187]=23504;
squeal_samples[11188]=25929;
squeal_samples[11189]=28251;
squeal_samples[11190]=30466;
squeal_samples[11191]=32593;
squeal_samples[11192]=34618;
squeal_samples[11193]=36559;
squeal_samples[11194]=38401;
squeal_samples[11195]=40174;
squeal_samples[11196]=41857;
squeal_samples[11197]=43476;
squeal_samples[11198]=45010;
squeal_samples[11199]=46488;
squeal_samples[11200]=47889;
squeal_samples[11201]=49235;
squeal_samples[11202]=50522;
squeal_samples[11203]=51747;
squeal_samples[11204]=52089;
squeal_samples[11205]=47523;
squeal_samples[11206]=42461;
squeal_samples[11207]=37711;
squeal_samples[11208]=33281;
squeal_samples[11209]=29121;
squeal_samples[11210]=25241;
squeal_samples[11211]=21601;
squeal_samples[11212]=18202;
squeal_samples[11213]=15020;
squeal_samples[11214]=12042;
squeal_samples[11215]=9256;
squeal_samples[11216]=6828;
squeal_samples[11217]=8412;
squeal_samples[11218]=11489;
squeal_samples[11219]=14437;
squeal_samples[11220]=17265;
squeal_samples[11221]=19966;
squeal_samples[11222]=22551;
squeal_samples[11223]=25023;
squeal_samples[11224]=27375;
squeal_samples[11225]=29636;
squeal_samples[11226]=31796;
squeal_samples[11227]=33855;
squeal_samples[11228]=35830;
squeal_samples[11229]=37703;
squeal_samples[11230]=39508;
squeal_samples[11231]=41221;
squeal_samples[11232]=42866;
squeal_samples[11233]=44431;
squeal_samples[11234]=45928;
squeal_samples[11235]=47356;
squeal_samples[11236]=48726;
squeal_samples[11237]=50028;
squeal_samples[11238]=51283;
squeal_samples[11239]=52419;
squeal_samples[11240]=49498;
squeal_samples[11241]=44305;
squeal_samples[11242]=39446;
squeal_samples[11243]=34891;
squeal_samples[11244]=30637;
squeal_samples[11245]=26647;
squeal_samples[11246]=22925;
squeal_samples[11247]=19436;
squeal_samples[11248]=16173;
squeal_samples[11249]=13121;
squeal_samples[11250]=10263;
squeal_samples[11251]=7591;
squeal_samples[11252]=7914;
squeal_samples[11253]=11011;
squeal_samples[11254]=13980;
squeal_samples[11255]=16825;
squeal_samples[11256]=19545;
squeal_samples[11257]=22148;
squeal_samples[11258]=24630;
squeal_samples[11259]=27008;
squeal_samples[11260]=29277;
squeal_samples[11261]=31455;
squeal_samples[11262]=33532;
squeal_samples[11263]=35510;
squeal_samples[11264]=37413;
squeal_samples[11265]=39220;
squeal_samples[11266]=40947;
squeal_samples[11267]=42604;
squeal_samples[11268]=44181;
squeal_samples[11269]=45687;
squeal_samples[11270]=47131;
squeal_samples[11271]=48503;
squeal_samples[11272]=49823;
squeal_samples[11273]=51072;
squeal_samples[11274]=52284;
squeal_samples[11275]=50889;
squeal_samples[11276]=45657;
squeal_samples[11277]=40708;
squeal_samples[11278]=36073;
squeal_samples[11279]=31739;
squeal_samples[11280]=27685;
squeal_samples[11281]=23891;
squeal_samples[11282]=20343;
squeal_samples[11283]=17016;
squeal_samples[11284]=13912;
squeal_samples[11285]=11004;
squeal_samples[11286]=8280;
squeal_samples[11287]=6846;
squeal_samples[11288]=9600;
squeal_samples[11289]=12631;
squeal_samples[11290]=15529;
squeal_samples[11291]=18306;
squeal_samples[11292]=20958;
squeal_samples[11293]=23503;
squeal_samples[11294]=25926;
squeal_samples[11295]=28246;
squeal_samples[11296]=30458;
squeal_samples[11297]=32583;
squeal_samples[11298]=34605;
squeal_samples[11299]=36543;
squeal_samples[11300]=38390;
squeal_samples[11301]=40154;
squeal_samples[11302]=41849;
squeal_samples[11303]=43456;
squeal_samples[11304]=44995;
squeal_samples[11305]=46464;
squeal_samples[11306]=47873;
squeal_samples[11307]=49213;
squeal_samples[11308]=50497;
squeal_samples[11309]=51723;
squeal_samples[11310]=52060;
squeal_samples[11311]=47504;
squeal_samples[11312]=42428;
squeal_samples[11313]=37694;
squeal_samples[11314]=33242;
squeal_samples[11315]=29096;
squeal_samples[11316]=25206;
squeal_samples[11317]=21574;
squeal_samples[11318]=18169;
squeal_samples[11319]=14985;
squeal_samples[11320]=12005;
squeal_samples[11321]=9223;
squeal_samples[11322]=7018;
squeal_samples[11323]=9067;
squeal_samples[11324]=12125;
squeal_samples[11325]=15033;
squeal_samples[11326]=17840;
squeal_samples[11327]=20507;
squeal_samples[11328]=23073;
squeal_samples[11329]=25513;
squeal_samples[11330]=27855;
squeal_samples[11331]=30079;
squeal_samples[11332]=32223;
squeal_samples[11333]=34259;
squeal_samples[11334]=36209;
squeal_samples[11335]=38077;
squeal_samples[11336]=39855;
squeal_samples[11337]=41556;
squeal_samples[11338]=43178;
squeal_samples[11339]=44728;
squeal_samples[11340]=46215;
squeal_samples[11341]=47627;
squeal_samples[11342]=48985;
squeal_samples[11343]=50271;
squeal_samples[11344]=51503;
squeal_samples[11345]=52486;
squeal_samples[11346]=48892;
squeal_samples[11347]=43741;
squeal_samples[11348]=38907;
squeal_samples[11349]=34390;
squeal_samples[11350]=30165;
squeal_samples[11351]=26211;
squeal_samples[11352]=22507;
squeal_samples[11353]=19044;
squeal_samples[11354]=15799;
squeal_samples[11355]=12772;
squeal_samples[11356]=9932;
squeal_samples[11357]=7284;
squeal_samples[11358]=7619;
squeal_samples[11359]=10725;
squeal_samples[11360]=13705;
squeal_samples[11361]=16557;
squeal_samples[11362]=19285;
squeal_samples[11363]=21902;
squeal_samples[11364]=24392;
squeal_samples[11365]=26784;
squeal_samples[11366]=29055;
squeal_samples[11367]=31242;
squeal_samples[11368]=33325;
squeal_samples[11369]=35314;
squeal_samples[11370]=37219;
squeal_samples[11371]=39031;
squeal_samples[11372]=40772;
squeal_samples[11373]=42430;
squeal_samples[11374]=44017;
squeal_samples[11375]=45531;
squeal_samples[11376]=46974;
squeal_samples[11377]=48357;
squeal_samples[11378]=49672;
squeal_samples[11379]=50940;
squeal_samples[11380]=52139;
squeal_samples[11381]=51425;
squeal_samples[11382]=46308;
squeal_samples[11383]=41307;
squeal_samples[11384]=36641;
squeal_samples[11385]=32259;
squeal_samples[11386]=28172;
squeal_samples[11387]=24343;
squeal_samples[11388]=20762;
squeal_samples[11389]=17410;
squeal_samples[11390]=14273;
squeal_samples[11391]=11337;
squeal_samples[11392]=8593;
squeal_samples[11393]=6738;
squeal_samples[11394]=9190;
squeal_samples[11395]=12235;
squeal_samples[11396]=15152;
squeal_samples[11397]=17943;
squeal_samples[11398]=20609;
squeal_samples[11399]=23161;
squeal_samples[11400]=25604;
squeal_samples[11401]=27931;
squeal_samples[11402]=30165;
squeal_samples[11403]=32294;
squeal_samples[11404]=34331;
squeal_samples[11405]=36275;
squeal_samples[11406]=38134;
squeal_samples[11407]=39910;
squeal_samples[11408]=41610;
squeal_samples[11409]=43224;
squeal_samples[11410]=44780;
squeal_samples[11411]=46255;
squeal_samples[11412]=47666;
squeal_samples[11413]=49017;
squeal_samples[11414]=50306;
squeal_samples[11415]=51540;
squeal_samples[11416]=52507;
squeal_samples[11417]=48923;
squeal_samples[11418]=43759;
squeal_samples[11419]=38930;
squeal_samples[11420]=34406;
squeal_samples[11421]=30174;
squeal_samples[11422]=26222;
squeal_samples[11423]=22512;
squeal_samples[11424]=19048;
squeal_samples[11425]=15806;
squeal_samples[11426]=12768;
squeal_samples[11427]=9934;
squeal_samples[11428]=7279;
squeal_samples[11429]=7609;
squeal_samples[11430]=10723;
squeal_samples[11431]=13696;
squeal_samples[11432]=16552;
squeal_samples[11433]=19281;
squeal_samples[11434]=21886;
squeal_samples[11435]=24386;
squeal_samples[11436]=26767;
squeal_samples[11437]=29048;
squeal_samples[11438]=31229;
squeal_samples[11439]=33312;
squeal_samples[11440]=35305;
squeal_samples[11441]=37205;
squeal_samples[11442]=39022;
squeal_samples[11443]=40759;
squeal_samples[11444]=42414;
squeal_samples[11445]=43999;
squeal_samples[11446]=45515;
squeal_samples[11447]=46957;
squeal_samples[11448]=48339;
squeal_samples[11449]=49657;
squeal_samples[11450]=50916;
squeal_samples[11451]=52123;
squeal_samples[11452]=51408;
squeal_samples[11453]=46285;
squeal_samples[11454]=41287;
squeal_samples[11455]=36621;
squeal_samples[11456]=32239;
squeal_samples[11457]=28153;
squeal_samples[11458]=24322;
squeal_samples[11459]=20740;
squeal_samples[11460]=17388;
squeal_samples[11461]=14250;
squeal_samples[11462]=11314;
squeal_samples[11463]=8572;
squeal_samples[11464]=6714;
squeal_samples[11465]=9171;
squeal_samples[11466]=12210;
squeal_samples[11467]=15131;
squeal_samples[11468]=17914;
squeal_samples[11469]=20588;
squeal_samples[11470]=23138;
squeal_samples[11471]=25581;
squeal_samples[11472]=27905;
squeal_samples[11473]=30135;
squeal_samples[11474]=32268;
squeal_samples[11475]=34303;
squeal_samples[11476]=36252;
squeal_samples[11477]=38107;
squeal_samples[11478]=39888;
squeal_samples[11479]=41580;
squeal_samples[11480]=43205;
squeal_samples[11481]=44750;
squeal_samples[11482]=46228;
squeal_samples[11483]=47640;
squeal_samples[11484]=48991;
squeal_samples[11485]=50281;
squeal_samples[11486]=51511;
squeal_samples[11487]=52480;
squeal_samples[11488]=48896;
squeal_samples[11489]=43729;
squeal_samples[11490]=38904;
squeal_samples[11491]=34376;
squeal_samples[11492]=30149;
squeal_samples[11493]=26193;
squeal_samples[11494]=22489;
squeal_samples[11495]=19022;
squeal_samples[11496]=15775;
squeal_samples[11497]=12744;
squeal_samples[11498]=9903;
squeal_samples[11499]=7254;
squeal_samples[11500]=7580;
squeal_samples[11501]=10695;
squeal_samples[11502]=13670;
squeal_samples[11503]=16521;
squeal_samples[11504]=19257;
squeal_samples[11505]=21861;
squeal_samples[11506]=24361;
squeal_samples[11507]=26736;
squeal_samples[11508]=29024;
squeal_samples[11509]=31197;
squeal_samples[11510]=33288;
squeal_samples[11511]=35276;
squeal_samples[11512]=37176;
squeal_samples[11513]=38996;
squeal_samples[11514]=40730;
squeal_samples[11515]=42387;
squeal_samples[11516]=43971;
squeal_samples[11517]=45487;
squeal_samples[11518]=46930;
squeal_samples[11519]=48310;
squeal_samples[11520]=49631;
squeal_samples[11521]=50892;
squeal_samples[11522]=52096;
squeal_samples[11523]=51381;
squeal_samples[11524]=46255;
squeal_samples[11525]=41261;
squeal_samples[11526]=36593;
squeal_samples[11527]=32210;
squeal_samples[11528]=28128;
squeal_samples[11529]=24291;
squeal_samples[11530]=20715;
squeal_samples[11531]=17358;
squeal_samples[11532]=14223;
squeal_samples[11533]=11287;
squeal_samples[11534]=8543;
squeal_samples[11535]=6687;
squeal_samples[11536]=9143;
squeal_samples[11537]=12182;
squeal_samples[11538]=15103;
squeal_samples[11539]=17887;
squeal_samples[11540]=20558;
squeal_samples[11541]=23113;
squeal_samples[11542]=25552;
squeal_samples[11543]=27882;
squeal_samples[11544]=30108;
squeal_samples[11545]=32239;
squeal_samples[11546]=34277;
squeal_samples[11547]=36222;
squeal_samples[11548]=38081;
squeal_samples[11549]=39858;
squeal_samples[11550]=41555;
squeal_samples[11551]=43174;
squeal_samples[11552]=44725;
squeal_samples[11553]=46197;
squeal_samples[11554]=47615;
squeal_samples[11555]=48961;
squeal_samples[11556]=50255;
squeal_samples[11557]=51482;
squeal_samples[11558]=52451;
squeal_samples[11559]=48871;
squeal_samples[11560]=43698;
squeal_samples[11561]=38880;
squeal_samples[11562]=34344;
squeal_samples[11563]=30123;
squeal_samples[11564]=26163;
squeal_samples[11565]=22464;
squeal_samples[11566]=18991;
squeal_samples[11567]=15750;
squeal_samples[11568]=12713;
squeal_samples[11569]=9876;
squeal_samples[11570]=7272;
squeal_samples[11571]=8255;
squeal_samples[11572]=11335;
squeal_samples[11573]=14282;
squeal_samples[11574]=17109;
squeal_samples[11575]=19810;
squeal_samples[11576]=22398;
squeal_samples[11577]=24865;
squeal_samples[11578]=27229;
squeal_samples[11579]=29484;
squeal_samples[11580]=31641;
squeal_samples[11581]=33702;
squeal_samples[11582]=35678;
squeal_samples[11583]=37555;
squeal_samples[11584]=39358;
squeal_samples[11585]=41071;
squeal_samples[11586]=42719;
squeal_samples[11587]=44283;
squeal_samples[11588]=45787;
squeal_samples[11589]=47208;
squeal_samples[11590]=48584;
squeal_samples[11591]=49883;
squeal_samples[11592]=51132;
squeal_samples[11593]=52323;
squeal_samples[11594]=50935;
squeal_samples[11595]=45682;
squeal_samples[11596]=40730;
squeal_samples[11597]=36084;
squeal_samples[11598]=31740;
squeal_samples[11599]=27679;
squeal_samples[11600]=23875;
squeal_samples[11601]=20321;
squeal_samples[11602]=16989;
squeal_samples[11603]=13873;
squeal_samples[11604]=10962;
squeal_samples[11605]=8237;
squeal_samples[11606]=6797;
squeal_samples[11607]=9546;
squeal_samples[11608]=12569;
squeal_samples[11609]=15472;
squeal_samples[11610]=18238;
squeal_samples[11611]=20898;
squeal_samples[11612]=23426;
squeal_samples[11613]=25861;
squeal_samples[11614]=28165;
squeal_samples[11615]=30387;
squeal_samples[11616]=32502;
squeal_samples[11617]=34527;
squeal_samples[11618]=36460;
squeal_samples[11619]=38308;
squeal_samples[11620]=40069;
squeal_samples[11621]=41760;
squeal_samples[11622]=43364;
squeal_samples[11623]=44908;
squeal_samples[11624]=46371;
squeal_samples[11625]=47782;
squeal_samples[11626]=49118;
squeal_samples[11627]=50402;
squeal_samples[11628]=51620;
squeal_samples[11629]=52331;
squeal_samples[11630]=48190;
squeal_samples[11631]=43073;
squeal_samples[11632]=38276;
squeal_samples[11633]=33794;
squeal_samples[11634]=29599;
squeal_samples[11635]=25669;
squeal_samples[11636]=21996;
squeal_samples[11637]=18555;
squeal_samples[11638]=15342;
squeal_samples[11639]=12333;
squeal_samples[11640]=9516;
squeal_samples[11641]=7065;
squeal_samples[11642]=8624;
squeal_samples[11643]=11692;
squeal_samples[11644]=14624;
squeal_samples[11645]=17434;
squeal_samples[11646]=20119;
squeal_samples[11647]=22691;
squeal_samples[11648]=25146;
squeal_samples[11649]=27494;
squeal_samples[11650]=29733;
squeal_samples[11651]=31884;
squeal_samples[11652]=33935;
squeal_samples[11653]=35895;
squeal_samples[11654]=37760;
squeal_samples[11655]=39552;
squeal_samples[11656]=41262;
squeal_samples[11657]=42888;
squeal_samples[11658]=44455;
squeal_samples[11659]=45939;
squeal_samples[11660]=47365;
squeal_samples[11661]=48719;
squeal_samples[11662]=50024;
squeal_samples[11663]=51256;
squeal_samples[11664]=52452;
squeal_samples[11665]=50274;
squeal_samples[11666]=45020;
squeal_samples[11667]=40105;
squeal_samples[11668]=35501;
squeal_samples[11669]=31192;
squeal_samples[11670]=27161;
squeal_samples[11671]=23391;
squeal_samples[11672]=19864;
squeal_samples[11673]=16560;
squeal_samples[11674]=13475;
squeal_samples[11675]=10588;
squeal_samples[11676]=7879;
squeal_samples[11677]=6946;
squeal_samples[11678]=9902;
squeal_samples[11679]=12919;
squeal_samples[11680]=15794;
squeal_samples[11681]=18554;
squeal_samples[11682]=21194;
squeal_samples[11683]=23710;
squeal_samples[11684]=26129;
squeal_samples[11685]=28422;
squeal_samples[11686]=30628;
squeal_samples[11687]=32731;
squeal_samples[11688]=34749;
squeal_samples[11689]=36663;
squeal_samples[11690]=38511;
squeal_samples[11691]=40256;
squeal_samples[11692]=41940;
squeal_samples[11693]=43535;
squeal_samples[11694]=45066;
squeal_samples[11695]=46523;
squeal_samples[11696]=47918;
squeal_samples[11697]=49258;
squeal_samples[11698]=50526;
squeal_samples[11699]=51750;
squeal_samples[11700]=52439;
squeal_samples[11701]=48295;
squeal_samples[11702]=43168;
squeal_samples[11703]=38368;
squeal_samples[11704]=33877;
squeal_samples[11705]=29670;
squeal_samples[11706]=25742;
squeal_samples[11707]=22059;
squeal_samples[11708]=18615;
squeal_samples[11709]=15390;
squeal_samples[11710]=12375;
squeal_samples[11711]=9560;
squeal_samples[11712]=6967;
squeal_samples[11713]=7961;
squeal_samples[11714]=11054;
squeal_samples[11715]=14016;
squeal_samples[11716]=16847;
squeal_samples[11717]=19559;
squeal_samples[11718]=22152;
squeal_samples[11719]=24630;
squeal_samples[11720]=26999;
squeal_samples[11721]=29261;
squeal_samples[11722]=31428;
squeal_samples[11723]=33497;
squeal_samples[11724]=35479;
squeal_samples[11725]=37360;
squeal_samples[11726]=39175;
squeal_samples[11727]=40890;
squeal_samples[11728]=42541;
squeal_samples[11729]=44116;
squeal_samples[11730]=45613;
squeal_samples[11731]=47054;
squeal_samples[11732]=48422;
squeal_samples[11733]=49730;
squeal_samples[11734]=50988;
squeal_samples[11735]=52180;
squeal_samples[11736]=51460;
squeal_samples[11737]=46323;
squeal_samples[11738]=41325;
squeal_samples[11739]=36636;
squeal_samples[11740]=32256;
squeal_samples[11741]=28152;
squeal_samples[11742]=24321;
squeal_samples[11743]=20730;
squeal_samples[11744]=17369;
squeal_samples[11745]=14231;
squeal_samples[11746]=11283;
squeal_samples[11747]=8542;
squeal_samples[11748]=6673;
squeal_samples[11749]=9129;
squeal_samples[11750]=12164;
squeal_samples[11751]=15079;
squeal_samples[11752]=17867;
squeal_samples[11753]=20537;
squeal_samples[11754]=23079;
squeal_samples[11755]=25525;
squeal_samples[11756]=27847;
squeal_samples[11757]=30072;
squeal_samples[11758]=32205;
squeal_samples[11759]=34240;
squeal_samples[11760]=36184;
squeal_samples[11761]=38037;
squeal_samples[11762]=39816;
squeal_samples[11763]=41505;
squeal_samples[11764]=43125;
squeal_samples[11765]=44672;
squeal_samples[11766]=46147;
squeal_samples[11767]=47561;
squeal_samples[11768]=48907;
squeal_samples[11769]=50195;
squeal_samples[11770]=51426;
squeal_samples[11771]=52553;
squeal_samples[11772]=49613;
squeal_samples[11773]=44398;
squeal_samples[11774]=39516;
squeal_samples[11775]=34952;
squeal_samples[11776]=30669;
squeal_samples[11777]=26674;
squeal_samples[11778]=22932;
squeal_samples[11779]=19430;
squeal_samples[11780]=16154;
squeal_samples[11781]=13085;
squeal_samples[11782]=10224;
squeal_samples[11783]=7540;
squeal_samples[11784]=7195;
squeal_samples[11785]=10270;
squeal_samples[11786]=13260;
squeal_samples[11787]=16128;
squeal_samples[11788]=18864;
squeal_samples[11789]=21488;
squeal_samples[11790]=23994;
squeal_samples[11791]=26390;
squeal_samples[11792]=28679;
squeal_samples[11793]=30873;
squeal_samples[11794]=32960;
squeal_samples[11795]=34966;
squeal_samples[11796]=36873;
squeal_samples[11797]=38698;
squeal_samples[11798]=40446;
squeal_samples[11799]=42110;
squeal_samples[11800]=43703;
squeal_samples[11801]=45223;
squeal_samples[11802]=46668;
squeal_samples[11803]=48066;
squeal_samples[11804]=49378;
squeal_samples[11805]=50652;
squeal_samples[11806]=51862;
squeal_samples[11807]=52186;
squeal_samples[11808]=47606;
squeal_samples[11809]=42512;
squeal_samples[11810]=37756;
squeal_samples[11811]=33295;
squeal_samples[11812]=29125;
squeal_samples[11813]=25231;
squeal_samples[11814]=21576;
squeal_samples[11815]=18162;
squeal_samples[11816]=14966;
squeal_samples[11817]=11975;
squeal_samples[11818]=9180;
squeal_samples[11819]=6745;
squeal_samples[11820]=8314;
squeal_samples[11821]=11396;
squeal_samples[11822]=14335;
squeal_samples[11823]=17157;
squeal_samples[11824]=19850;
squeal_samples[11825]=22427;
squeal_samples[11826]=24894;
squeal_samples[11827]=27250;
squeal_samples[11828]=29499;
squeal_samples[11829]=31652;
squeal_samples[11830]=33712;
squeal_samples[11831]=35676;
squeal_samples[11832]=37556;
squeal_samples[11833]=39351;
squeal_samples[11834]=41061;
squeal_samples[11835]=42700;
squeal_samples[11836]=44262;
squeal_samples[11837]=45757;
squeal_samples[11838]=47183;
squeal_samples[11839]=48550;
squeal_samples[11840]=49849;
squeal_samples[11841]=51099;
squeal_samples[11842]=52290;
squeal_samples[11843]=50890;
squeal_samples[11844]=45640;
squeal_samples[11845]=40678;
squeal_samples[11846]=36036;
squeal_samples[11847]=31684;
squeal_samples[11848]=27619;
squeal_samples[11849]=23814;
squeal_samples[11850]=20254;
squeal_samples[11851]=16925;
squeal_samples[11852]=13805;
squeal_samples[11853]=10893;
squeal_samples[11854]=8162;
squeal_samples[11855]=6723;
squeal_samples[11856]=9467;
squeal_samples[11857]=12500;
squeal_samples[11858]=15392;
squeal_samples[11859]=18165;
squeal_samples[11860]=20816;
squeal_samples[11861]=23356;
squeal_samples[11862]=25770;
squeal_samples[11863]=28090;
squeal_samples[11864]=30305;
squeal_samples[11865]=32424;
squeal_samples[11866]=34442;
squeal_samples[11867]=36373;
squeal_samples[11868]=38224;
squeal_samples[11869]=39989;
squeal_samples[11870]=41670;
squeal_samples[11871]=43283;
squeal_samples[11872]=44818;
squeal_samples[11873]=46286;
squeal_samples[11874]=47689;
squeal_samples[11875]=49030;
squeal_samples[11876]=50308;
squeal_samples[11877]=51536;
squeal_samples[11878]=52495;
squeal_samples[11879]=48896;
squeal_samples[11880]=43729;
squeal_samples[11881]=38888;
squeal_samples[11882]=34354;
squeal_samples[11883]=30117;
squeal_samples[11884]=26147;
squeal_samples[11885]=22439;
squeal_samples[11886]=18966;
squeal_samples[11887]=15719;
squeal_samples[11888]=12674;
squeal_samples[11889]=9836;
squeal_samples[11890]=7216;
squeal_samples[11891]=8203;
squeal_samples[11892]=11275;
squeal_samples[11893]=14228;
squeal_samples[11894]=17045;
squeal_samples[11895]=19746;
squeal_samples[11896]=22328;
squeal_samples[11897]=24800;
squeal_samples[11898]=27148;
squeal_samples[11899]=29409;
squeal_samples[11900]=31560;
squeal_samples[11901]=33627;
squeal_samples[11902]=35591;
squeal_samples[11903]=37474;
squeal_samples[11904]=39267;
squeal_samples[11905]=40989;
squeal_samples[11906]=42629;
squeal_samples[11907]=44189;
squeal_samples[11908]=45691;
squeal_samples[11909]=47116;
squeal_samples[11910]=48481;
squeal_samples[11911]=49785;
squeal_samples[11912]=51035;
squeal_samples[11913]=52224;
squeal_samples[11914]=51497;
squeal_samples[11915]=46355;
squeal_samples[11916]=41345;
squeal_samples[11917]=36659;
squeal_samples[11918]=32269;
squeal_samples[11919]=28160;
squeal_samples[11920]=24323;
squeal_samples[11921]=20726;
squeal_samples[11922]=17362;
squeal_samples[11923]=14219;
squeal_samples[11924]=11272;
squeal_samples[11925]=8520;
squeal_samples[11926]=6650;
squeal_samples[11927]=9108;
squeal_samples[11928]=12139;
squeal_samples[11929]=15053;
squeal_samples[11930]=17833;
squeal_samples[11931]=20503;
squeal_samples[11932]=23048;
squeal_samples[11933]=25483;
squeal_samples[11934]=27811;
squeal_samples[11935]=30036;
squeal_samples[11936]=32169;
squeal_samples[11937]=34194;
squeal_samples[11938]=36140;
squeal_samples[11939]=37994;
squeal_samples[11940]=39770;
squeal_samples[11941]=41463;
squeal_samples[11942]=43079;
squeal_samples[11943]=44624;
squeal_samples[11944]=46095;
squeal_samples[11945]=47515;
squeal_samples[11946]=48853;
squeal_samples[11947]=50150;
squeal_samples[11948]=51372;
squeal_samples[11949]=52500;
squeal_samples[11950]=49558;
squeal_samples[11951]=44341;
squeal_samples[11952]=39458;
squeal_samples[11953]=34890;
squeal_samples[11954]=30614;
squeal_samples[11955]=26614;
squeal_samples[11956]=22869;
squeal_samples[11957]=19371;
squeal_samples[11958]=16093;
squeal_samples[11959]=13024;
squeal_samples[11960]=10157;
squeal_samples[11961]=7473;
squeal_samples[11962]=7786;
squeal_samples[11963]=10879;
squeal_samples[11964]=13838;
squeal_samples[11965]=16683;
squeal_samples[11966]=19387;
squeal_samples[11967]=21994;
squeal_samples[11968]=24470;
squeal_samples[11969]=26839;
squeal_samples[11970]=29109;
squeal_samples[11971]=31275;
squeal_samples[11972]=33349;
squeal_samples[11973]=35324;
squeal_samples[11974]=37223;
squeal_samples[11975]=39026;
squeal_samples[11976]=40755;
squeal_samples[11977]=42397;
squeal_samples[11978]=43980;
squeal_samples[11979]=45478;
squeal_samples[11980]=46919;
squeal_samples[11981]=48285;
squeal_samples[11982]=49601;
squeal_samples[11983]=50854;
squeal_samples[11984]=52052;
squeal_samples[11985]=51899;
squeal_samples[11986]=46978;
squeal_samples[11987]=41925;
squeal_samples[11988]=37201;
squeal_samples[11989]=32772;
squeal_samples[11990]=28635;
squeal_samples[11991]=24765;
squeal_samples[11992]=21132;
squeal_samples[11993]=17747;
squeal_samples[11994]=14563;
squeal_samples[11995]=11610;
squeal_samples[11996]=8821;
squeal_samples[11997]=6632;
squeal_samples[11998]=8684;
squeal_samples[11999]=11738;
squeal_samples[12000]=14670;
squeal_samples[12001]=17463;
squeal_samples[12002]=20148;
squeal_samples[12003]=22709;
squeal_samples[12004]=25157;
squeal_samples[12005]=27499;
squeal_samples[12006]=29732;
squeal_samples[12007]=31879;
squeal_samples[12008]=33915;
squeal_samples[12009]=35873;
squeal_samples[12010]=37737;
squeal_samples[12011]=39525;
squeal_samples[12012]=41227;
squeal_samples[12013]=42851;
squeal_samples[12014]=44407;
squeal_samples[12015]=45892;
squeal_samples[12016]=47306;
squeal_samples[12017]=48667;
squeal_samples[12018]=49958;
squeal_samples[12019]=51195;
squeal_samples[12020]=52373;
squeal_samples[12021]=50974;
squeal_samples[12022]=45711;
squeal_samples[12023]=40746;
squeal_samples[12024]=36085;
squeal_samples[12025]=31734;
squeal_samples[12026]=27659;
squeal_samples[12027]=23847;
squeal_samples[12028]=20281;
squeal_samples[12029]=16942;
squeal_samples[12030]=13825;
squeal_samples[12031]=10896;
squeal_samples[12032]=8173;
squeal_samples[12033]=6715;
squeal_samples[12034]=9471;
squeal_samples[12035]=12490;
squeal_samples[12036]=15381;
squeal_samples[12037]=18152;
squeal_samples[12038]=20798;
squeal_samples[12039]=23339;
squeal_samples[12040]=25752;
squeal_samples[12041]=28068;
squeal_samples[12042]=30275;
squeal_samples[12043]=32396;
squeal_samples[12044]=34413;
squeal_samples[12045]=36344;
squeal_samples[12046]=38192;
squeal_samples[12047]=39953;
squeal_samples[12048]=41637;
squeal_samples[12049]=43243;
squeal_samples[12050]=44779;
squeal_samples[12051]=46245;
squeal_samples[12052]=47647;
squeal_samples[12053]=48986;
squeal_samples[12054]=50267;
squeal_samples[12055]=51489;
squeal_samples[12056]=52606;
squeal_samples[12057]=49658;
squeal_samples[12058]=44427;
squeal_samples[12059]=39539;
squeal_samples[12060]=34967;
squeal_samples[12061]=30678;
squeal_samples[12062]=26674;
squeal_samples[12063]=22926;
squeal_samples[12064]=19417;
squeal_samples[12065]=16133;
squeal_samples[12066]=13057;
squeal_samples[12067]=10188;
squeal_samples[12068]=7504;
squeal_samples[12069]=7148;
squeal_samples[12070]=10222;
squeal_samples[12071]=13210;
squeal_samples[12072]=16072;
squeal_samples[12073]=18815;
squeal_samples[12074]=21432;
squeal_samples[12075]=23934;
squeal_samples[12076]=26329;
squeal_samples[12077]=28612;
squeal_samples[12078]=30808;
squeal_samples[12079]=32892;
squeal_samples[12080]=34897;
squeal_samples[12081]=36798;
squeal_samples[12082]=38630;
squeal_samples[12083]=40366;
squeal_samples[12084]=42029;
squeal_samples[12085]=43621;
squeal_samples[12086]=45137;
squeal_samples[12087]=46591;
squeal_samples[12088]=47971;
squeal_samples[12089]=49302;
squeal_samples[12090]=50559;
squeal_samples[12091]=51775;
squeal_samples[12092]=52457;
squeal_samples[12093]=48304;
squeal_samples[12094]=43165;
squeal_samples[12095]=38355;
squeal_samples[12096]=33855;
squeal_samples[12097]=29638;
squeal_samples[12098]=25703;
squeal_samples[12099]=22010;
squeal_samples[12100]=18561;
squeal_samples[12101]=15329;
squeal_samples[12102]=12311;
squeal_samples[12103]=9481;
squeal_samples[12104]=6893;
squeal_samples[12105]=7878;
squeal_samples[12106]=10968;
squeal_samples[12107]=13923;
squeal_samples[12108]=16753;
squeal_samples[12109]=19462;
squeal_samples[12110]=22054;
squeal_samples[12111]=24532;
squeal_samples[12112]=26896;
squeal_samples[12113]=29156;
squeal_samples[12114]=31324;
squeal_samples[12115]=33391;
squeal_samples[12116]=35366;
squeal_samples[12117]=37250;
squeal_samples[12118]=39050;
squeal_samples[12119]=40778;
squeal_samples[12120]=42420;
squeal_samples[12121]=43992;
squeal_samples[12122]=45491;
squeal_samples[12123]=46929;
squeal_samples[12124]=48295;
squeal_samples[12125]=49606;
squeal_samples[12126]=50855;
squeal_samples[12127]=52055;
squeal_samples[12128]=51892;
squeal_samples[12129]=46972;
squeal_samples[12130]=41913;
squeal_samples[12131]=37186;
squeal_samples[12132]=32758;
squeal_samples[12133]=28615;
squeal_samples[12134]=24743;
squeal_samples[12135]=21109;
squeal_samples[12136]=17715;
squeal_samples[12137]=14545;
squeal_samples[12138]=11572;
squeal_samples[12139]=8795;
squeal_samples[12140]=6598;
squeal_samples[12141]=8651;
squeal_samples[12142]=11706;
squeal_samples[12143]=14628;
squeal_samples[12144]=17431;
squeal_samples[12145]=20108;
squeal_samples[12146]=22669;
squeal_samples[12147]=25119;
squeal_samples[12148]=27457;
squeal_samples[12149]=29689;
squeal_samples[12150]=31837;
squeal_samples[12151]=33874;
squeal_samples[12152]=35830;
squeal_samples[12153]=37695;
squeal_samples[12154]=39477;
squeal_samples[12155]=41178;
squeal_samples[12156]=42805;
squeal_samples[12157]=44359;
squeal_samples[12158]=45844;
squeal_samples[12159]=47259;
squeal_samples[12160]=48613;
squeal_samples[12161]=49904;
squeal_samples[12162]=51148;
squeal_samples[12163]=52328;
squeal_samples[12164]=50921;
squeal_samples[12165]=45663;
squeal_samples[12166]=40686;
squeal_samples[12167]=36038;
squeal_samples[12168]=31677;
squeal_samples[12169]=27608;
squeal_samples[12170]=23791;
squeal_samples[12171]=20229;
squeal_samples[12172]=16882;
squeal_samples[12173]=13767;
squeal_samples[12174]=10842;
squeal_samples[12175]=8112;
squeal_samples[12176]=7148;
squeal_samples[12177]=10093;
squeal_samples[12178]=13087;
squeal_samples[12179]=15949;
squeal_samples[12180]=18697;
squeal_samples[12181]=21315;
squeal_samples[12182]=23826;
squeal_samples[12183]=26219;
squeal_samples[12184]=28509;
squeal_samples[12185]=30702;
squeal_samples[12186]=32792;
squeal_samples[12187]=34794;
squeal_samples[12188]=36704;
squeal_samples[12189]=38534;
squeal_samples[12190]=40274;
squeal_samples[12191]=41942;
squeal_samples[12192]=43532;
squeal_samples[12193]=45051;
squeal_samples[12194]=46508;
squeal_samples[12195]=47891;
squeal_samples[12196]=49216;
squeal_samples[12197]=50486;
squeal_samples[12198]=51695;
squeal_samples[12199]=52382;
squeal_samples[12200]=48228;
squeal_samples[12201]=43091;
squeal_samples[12202]=38287;
squeal_samples[12203]=33781;
squeal_samples[12204]=29574;
squeal_samples[12205]=25636;
squeal_samples[12206]=21948;
squeal_samples[12207]=18498;
squeal_samples[12208]=15265;
squeal_samples[12209]=12254;
squeal_samples[12210]=9418;
squeal_samples[12211]=6967;
squeal_samples[12212]=8519;
squeal_samples[12213]=11576;
squeal_samples[12214]=14508;
squeal_samples[12215]=17312;
squeal_samples[12216]=19993;
squeal_samples[12217]=22557;
squeal_samples[12218]=25011;
squeal_samples[12219]=27348;
squeal_samples[12220]=29591;
squeal_samples[12221]=31736;
squeal_samples[12222]=33779;
squeal_samples[12223]=35738;
squeal_samples[12224]=37602;
squeal_samples[12225]=39396;
squeal_samples[12226]=41093;
squeal_samples[12227]=42728;
squeal_samples[12228]=44279;
squeal_samples[12229]=45768;
squeal_samples[12230]=47182;
squeal_samples[12231]=48544;
squeal_samples[12232]=49835;
squeal_samples[12233]=51081;
squeal_samples[12234]=52257;
squeal_samples[12235]=51526;
squeal_samples[12236]=46368;
squeal_samples[12237]=41353;
squeal_samples[12238]=36655;
squeal_samples[12239]=32258;
squeal_samples[12240]=28142;
squeal_samples[12241]=24296;
squeal_samples[12242]=20698;
squeal_samples[12243]=17321;
squeal_samples[12244]=14176;
squeal_samples[12245]=11222;
squeal_samples[12246]=8463;
squeal_samples[12247]=6592;
squeal_samples[12248]=9038;
squeal_samples[12249]=12078;
squeal_samples[12250]=14982;
squeal_samples[12251]=17764;
squeal_samples[12252]=20425;
squeal_samples[12253]=22970;
squeal_samples[12254]=25409;
squeal_samples[12255]=27731;
squeal_samples[12256]=29950;
squeal_samples[12257]=32079;
squeal_samples[12258]=34108;
squeal_samples[12259]=36050;
squeal_samples[12260]=37903;
squeal_samples[12261]=39674;
squeal_samples[12262]=41365;
squeal_samples[12263]=42980;
squeal_samples[12264]=44524;
squeal_samples[12265]=45998;
squeal_samples[12266]=47407;
squeal_samples[12267]=48751;
squeal_samples[12268]=50043;
squeal_samples[12269]=51269;
squeal_samples[12270]=52442;
squeal_samples[12271]=50265;
squeal_samples[12272]=44990;
squeal_samples[12273]=40060;
squeal_samples[12274]=35441;
squeal_samples[12275]=31124;
squeal_samples[12276]=27079;
squeal_samples[12277]=23305;
squeal_samples[12278]=19762;
squeal_samples[12279]=16451;
squeal_samples[12280]=13355;
squeal_samples[12281]=10457;
squeal_samples[12282]=7749;
squeal_samples[12283]=7371;
squeal_samples[12284]=10441;
squeal_samples[12285]=13411;
squeal_samples[12286]=16263;
squeal_samples[12287]=18985;
squeal_samples[12288]=21600;
squeal_samples[12289]=24090;
squeal_samples[12290]=26468;
squeal_samples[12291]=28747;
squeal_samples[12292]=30928;
squeal_samples[12293]=33009;
squeal_samples[12294]=34999;
squeal_samples[12295]=36899;
squeal_samples[12296]=38712;
squeal_samples[12297]=40446;
squeal_samples[12298]=42106;
squeal_samples[12299]=43680;
squeal_samples[12300]=45200;
squeal_samples[12301]=46638;
squeal_samples[12302]=48024;
squeal_samples[12303]=49333;
squeal_samples[12304]=50600;
squeal_samples[12305]=51796;
squeal_samples[12306]=52486;
squeal_samples[12307]=48316;
squeal_samples[12308]=43175;
squeal_samples[12309]=38354;
squeal_samples[12310]=33846;
squeal_samples[12311]=29633;
squeal_samples[12312]=25690;
squeal_samples[12313]=21990;
squeal_samples[12314]=18540;
squeal_samples[12315]=15299;
squeal_samples[12316]=12282;
squeal_samples[12317]=9449;
squeal_samples[12318]=6849;
squeal_samples[12319]=7842;
squeal_samples[12320]=10925;
squeal_samples[12321]=13882;
squeal_samples[12322]=16704;
squeal_samples[12323]=19420;
squeal_samples[12324]=22000;
squeal_samples[12325]=24478;
squeal_samples[12326]=26839;
squeal_samples[12327]=29101;
squeal_samples[12328]=31267;
squeal_samples[12329]=33329;
squeal_samples[12330]=35306;
squeal_samples[12331]=37186;
squeal_samples[12332]=38992;
squeal_samples[12333]=40707;
squeal_samples[12334]=42356;
squeal_samples[12335]=43928;
squeal_samples[12336]=45426;
squeal_samples[12337]=46861;
squeal_samples[12338]=48228;
squeal_samples[12339]=49539;
squeal_samples[12340]=50781;
squeal_samples[12341]=51983;
squeal_samples[12342]=52286;
squeal_samples[12343]=47687;
squeal_samples[12344]=42575;
squeal_samples[12345]=37803;
squeal_samples[12346]=33326;
squeal_samples[12347]=29139;
squeal_samples[12348]=25230;
squeal_samples[12349]=21564;
squeal_samples[12350]=18131;
squeal_samples[12351]=14924;
squeal_samples[12352]=11921;
squeal_samples[12353]=9121;
squeal_samples[12354]=6670;
squeal_samples[12355]=8239;
squeal_samples[12356]=11304;
squeal_samples[12357]=14244;
squeal_samples[12358]=17055;
squeal_samples[12359]=19746;
squeal_samples[12360]=22316;
squeal_samples[12361]=24785;
squeal_samples[12362]=27125;
squeal_samples[12363]=29382;
squeal_samples[12364]=31527;
squeal_samples[12365]=33582;
squeal_samples[12366]=35538;
squeal_samples[12367]=37418;
squeal_samples[12368]=39208;
squeal_samples[12369]=40916;
squeal_samples[12370]=42553;
squeal_samples[12371]=44113;
squeal_samples[12372]=45602;
squeal_samples[12373]=47030;
squeal_samples[12374]=48386;
squeal_samples[12375]=49689;
squeal_samples[12376]=50928;
squeal_samples[12377]=52122;
squeal_samples[12378]=51950;
squeal_samples[12379]=47019;
squeal_samples[12380]=41953;
squeal_samples[12381]=37216;
squeal_samples[12382]=32781;
squeal_samples[12383]=28624;
squeal_samples[12384]=24747;
squeal_samples[12385]=21109;
squeal_samples[12386]=17710;
squeal_samples[12387]=14527;
squeal_samples[12388]=11551;
squeal_samples[12389]=8764;
squeal_samples[12390]=6567;
squeal_samples[12391]=8612;
squeal_samples[12392]=11673;
squeal_samples[12393]=14589;
squeal_samples[12394]=17392;
squeal_samples[12395]=20058;
squeal_samples[12396]=22626;
squeal_samples[12397]=25069;
squeal_samples[12398]=27402;
squeal_samples[12399]=29634;
squeal_samples[12400]=31777;
squeal_samples[12401]=33813;
squeal_samples[12402]=35770;
squeal_samples[12403]=37629;
squeal_samples[12404]=39411;
squeal_samples[12405]=41112;
squeal_samples[12406]=42740;
squeal_samples[12407]=44286;
squeal_samples[12408]=45775;
squeal_samples[12409]=47185;
squeal_samples[12410]=48543;
squeal_samples[12411]=49834;
squeal_samples[12412]=51068;
squeal_samples[12413]=52251;
squeal_samples[12414]=51509;
squeal_samples[12415]=46354;
squeal_samples[12416]=41332;
squeal_samples[12417]=36630;
squeal_samples[12418]=32233;
squeal_samples[12419]=28109;
squeal_samples[12420]=24267;
squeal_samples[12421]=20658;
squeal_samples[12422]=17289;
squeal_samples[12423]=14131;
squeal_samples[12424]=11176;
squeal_samples[12425]=8422;
squeal_samples[12426]=6541;
squeal_samples[12427]=8994;
squeal_samples[12428]=12022;
squeal_samples[12429]=14932;
squeal_samples[12430]=17710;
squeal_samples[12431]=20371;
squeal_samples[12432]=22919;
squeal_samples[12433]=25354;
squeal_samples[12434]=27673;
squeal_samples[12435]=29898;
squeal_samples[12436]=32020;
squeal_samples[12437]=34050;
squeal_samples[12438]=35992;
squeal_samples[12439]=37842;
squeal_samples[12440]=39614;
squeal_samples[12441]=41303;
squeal_samples[12442]=42927;
squeal_samples[12443]=44459;
squeal_samples[12444]=45939;
squeal_samples[12445]=47345;
squeal_samples[12446]=48689;
squeal_samples[12447]=49979;
squeal_samples[12448]=51204;
squeal_samples[12449]=52378;
squeal_samples[12450]=50962;
squeal_samples[12451]=45691;
squeal_samples[12452]=40715;
squeal_samples[12453]=36050;
squeal_samples[12454]=31685;
squeal_samples[12455]=27601;
squeal_samples[12456]=23784;
squeal_samples[12457]=20210;
squeal_samples[12458]=16865;
squeal_samples[12459]=13737;
squeal_samples[12460]=10806;
squeal_samples[12461]=8071;
squeal_samples[12462]=6613;
squeal_samples[12463]=9365;
squeal_samples[12464]=12376;
squeal_samples[12465]=15270;
squeal_samples[12466]=18037;
squeal_samples[12467]=20682;
squeal_samples[12468]=23213;
squeal_samples[12469]=25632;
squeal_samples[12470]=27941;
squeal_samples[12471]=30153;
squeal_samples[12472]=32267;
squeal_samples[12473]=34281;
squeal_samples[12474]=36215;
squeal_samples[12475]=38051;
squeal_samples[12476]=39819;
squeal_samples[12477]=41493;
squeal_samples[12478]=43104;
squeal_samples[12479]=44634;
squeal_samples[12480]=46099;
squeal_samples[12481]=47500;
squeal_samples[12482]=48839;
squeal_samples[12483]=50111;
squeal_samples[12484]=51341;
squeal_samples[12485]=52501;
squeal_samples[12486]=50318;
squeal_samples[12487]=45035;
squeal_samples[12488]=40096;
squeal_samples[12489]=35469;
squeal_samples[12490]=31146;
squeal_samples[12491]=27093;
squeal_samples[12492]=23316;
squeal_samples[12493]=19762;
squeal_samples[12494]=16451;
squeal_samples[12495]=13339;
squeal_samples[12496]=10440;
squeal_samples[12497]=7725;
squeal_samples[12498]=7351;
squeal_samples[12499]=10407;
squeal_samples[12500]=13384;
squeal_samples[12501]=16231;
squeal_samples[12502]=18951;
squeal_samples[12503]=21557;
squeal_samples[12504]=24051;
squeal_samples[12505]=26423;
squeal_samples[12506]=28710;
squeal_samples[12507]=30880;
squeal_samples[12508]=32962;
squeal_samples[12509]=34949;
squeal_samples[12510]=36844;
squeal_samples[12511]=38662;
squeal_samples[12512]=40388;
squeal_samples[12513]=42049;
squeal_samples[12514]=43622;
squeal_samples[12515]=45142;
squeal_samples[12516]=46578;
squeal_samples[12517]=47958;
squeal_samples[12518]=49274;
squeal_samples[12519]=50532;
squeal_samples[12520]=51738;
squeal_samples[12521]=52414;
squeal_samples[12522]=48251;
squeal_samples[12523]=43106;
squeal_samples[12524]=38284;
squeal_samples[12525]=33780;
squeal_samples[12526]=29558;
squeal_samples[12527]=25609;
squeal_samples[12528]=21921;
squeal_samples[12529]=18455;
squeal_samples[12530]=15230;
squeal_samples[12531]=12199;
squeal_samples[12532]=9370;
squeal_samples[12533]=6902;
squeal_samples[12534]=8454;
squeal_samples[12535]=11514;
squeal_samples[12536]=14437;
squeal_samples[12537]=17238;
squeal_samples[12538]=19919;
squeal_samples[12539]=22481;
squeal_samples[12540]=24931;
squeal_samples[12541]=27268;
squeal_samples[12542]=29506;
squeal_samples[12543]=31649;
squeal_samples[12544]=33697;
squeal_samples[12545]=35646;
squeal_samples[12546]=37513;
squeal_samples[12547]=39292;
squeal_samples[12548]=41004;
squeal_samples[12549]=42625;
squeal_samples[12550]=44183;
squeal_samples[12551]=45659;
squeal_samples[12552]=47089;
squeal_samples[12553]=48433;
squeal_samples[12554]=49736;
squeal_samples[12555]=50966;
squeal_samples[12556]=52155;
squeal_samples[12557]=51415;
squeal_samples[12558]=46263;
squeal_samples[12559]=41244;
squeal_samples[12560]=36537;
squeal_samples[12561]=32146;
squeal_samples[12562]=28027;
squeal_samples[12563]=24179;
squeal_samples[12564]=20579;
squeal_samples[12565]=17203;
squeal_samples[12566]=14052;
squeal_samples[12567]=11097;
squeal_samples[12568]=8340;
squeal_samples[12569]=6869;
squeal_samples[12570]=9599;
squeal_samples[12571]=12605;
squeal_samples[12572]=15483;
squeal_samples[12573]=18245;
squeal_samples[12574]=20873;
squeal_samples[12575]=23399;
squeal_samples[12576]=25801;
squeal_samples[12577]=28110;
squeal_samples[12578]=30301;
squeal_samples[12579]=32414;
squeal_samples[12580]=34416;
squeal_samples[12581]=36342;
squeal_samples[12582]=38171;
squeal_samples[12583]=39928;
squeal_samples[12584]=41601;
squeal_samples[12585]=43203;
squeal_samples[12586]=44727;
squeal_samples[12587]=46192;
squeal_samples[12588]=47580;
squeal_samples[12589]=48909;
squeal_samples[12590]=50193;
squeal_samples[12591]=51397;
squeal_samples[12592]=52571;
squeal_samples[12593]=50366;
squeal_samples[12594]=45086;
squeal_samples[12595]=40136;
squeal_samples[12596]=35507;
squeal_samples[12597]=31176;
squeal_samples[12598]=27120;
squeal_samples[12599]=23336;
squeal_samples[12600]=19778;
squeal_samples[12601]=16459;
squeal_samples[12602]=13351;
squeal_samples[12603]=10447;
squeal_samples[12604]=7734;
squeal_samples[12605]=6775;
squeal_samples[12606]=9735;
squeal_samples[12607]=12729;
squeal_samples[12608]=15607;
squeal_samples[12609]=18351;
squeal_samples[12610]=20982;
squeal_samples[12611]=23498;
squeal_samples[12612]=25901;
squeal_samples[12613]=28192;
squeal_samples[12614]=30396;
squeal_samples[12615]=32490;
squeal_samples[12616]=34498;
squeal_samples[12617]=36410;
squeal_samples[12618]=38246;
squeal_samples[12619]=39993;
squeal_samples[12620]=41664;
squeal_samples[12621]=43261;
squeal_samples[12622]=44784;
squeal_samples[12623]=46243;
squeal_samples[12624]=47628;
squeal_samples[12625]=48964;
squeal_samples[12626]=50226;
squeal_samples[12627]=51442;
squeal_samples[12628]=52554;
squeal_samples[12629]=49591;
squeal_samples[12630]=44354;
squeal_samples[12631]=39452;
squeal_samples[12632]=34869;
squeal_samples[12633]=30572;
squeal_samples[12634]=26559;
squeal_samples[12635]=22803;
squeal_samples[12636]=19286;
squeal_samples[12637]=15999;
squeal_samples[12638]=12914;
squeal_samples[12639]=10040;
squeal_samples[12640]=7343;
squeal_samples[12641]=7646;
squeal_samples[12642]=10731;
squeal_samples[12643]=13695;
squeal_samples[12644]=16523;
squeal_samples[12645]=19235;
squeal_samples[12646]=21822;
squeal_samples[12647]=24299;
squeal_samples[12648]=26666;
squeal_samples[12649]=28927;
squeal_samples[12650]=31091;
squeal_samples[12651]=33155;
squeal_samples[12652]=35132;
squeal_samples[12653]=37020;
squeal_samples[12654]=38822;
squeal_samples[12655]=40548;
squeal_samples[12656]=42192;
squeal_samples[12657]=43761;
squeal_samples[12658]=45263;
squeal_samples[12659]=46700;
squeal_samples[12660]=48064;
squeal_samples[12661]=49379;
squeal_samples[12662]=50621;
squeal_samples[12663]=51829;
squeal_samples[12664]=52491;
squeal_samples[12665]=48330;
squeal_samples[12666]=43168;
squeal_samples[12667]=38340;
squeal_samples[12668]=33827;
squeal_samples[12669]=29602;
squeal_samples[12670]=25648;
squeal_samples[12671]=21945;
squeal_samples[12672]=18485;
squeal_samples[12673]=15242;
squeal_samples[12674]=12214;
squeal_samples[12675]=9377;
squeal_samples[12676]=6911;
squeal_samples[12677]=8450;
squeal_samples[12678]=11516;
squeal_samples[12679]=14431;
squeal_samples[12680]=17232;
squeal_samples[12681]=19908;
squeal_samples[12682]=22471;
squeal_samples[12683]=24918;
squeal_samples[12684]=27254;
squeal_samples[12685]=29488;
squeal_samples[12686]=31627;
squeal_samples[12687]=33675;
squeal_samples[12688]=35620;
squeal_samples[12689]=37489;
squeal_samples[12690]=39268;
squeal_samples[12691]=40972;
squeal_samples[12692]=42596;
squeal_samples[12693]=44147;
squeal_samples[12694]=45636;
squeal_samples[12695]=47050;
squeal_samples[12696]=48406;
squeal_samples[12697]=49697;
squeal_samples[12698]=50932;
squeal_samples[12699]=52114;
squeal_samples[12700]=51943;
squeal_samples[12701]=47000;
squeal_samples[12702]=41930;
squeal_samples[12703]=37181;
squeal_samples[12704]=32740;
squeal_samples[12705]=28580;
squeal_samples[12706]=24694;
squeal_samples[12707]=21057;
squeal_samples[12708]=17643;
squeal_samples[12709]=14464;
squeal_samples[12710]=11479;
squeal_samples[12711]=8691;
squeal_samples[12712]=6794;
squeal_samples[12713]=9223;
squeal_samples[12714]=12247;
squeal_samples[12715]=15135;
squeal_samples[12716]=17908;
squeal_samples[12717]=20547;
squeal_samples[12718]=23088;
squeal_samples[12719]=25499;
squeal_samples[12720]=27815;
squeal_samples[12721]=30022;
squeal_samples[12722]=32139;
squeal_samples[12723]=34157;
squeal_samples[12724]=36084;
squeal_samples[12725]=37930;
squeal_samples[12726]=39692;
squeal_samples[12727]=41378;
squeal_samples[12728]=42979;
squeal_samples[12729]=44514;
squeal_samples[12730]=45984;
squeal_samples[12731]=47378;
squeal_samples[12732]=48724;
squeal_samples[12733]=49995;
squeal_samples[12734]=51224;
squeal_samples[12735]=52386;
squeal_samples[12736]=50968;
squeal_samples[12737]=45687;
squeal_samples[12738]=40700;
squeal_samples[12739]=36032;
squeal_samples[12740]=31658;
squeal_samples[12741]=27574;
squeal_samples[12742]=23745;
squeal_samples[12743]=20169;
squeal_samples[12744]=16816;
squeal_samples[12745]=13679;
squeal_samples[12746]=10756;
squeal_samples[12747]=8005;
squeal_samples[12748]=7041;
squeal_samples[12749]=9975;
squeal_samples[12750]=12965;
squeal_samples[12751]=15827;
squeal_samples[12752]=18564;
squeal_samples[12753]=21182;
squeal_samples[12754]=23684;
squeal_samples[12755]=26072;
squeal_samples[12756]=28364;
squeal_samples[12757]=30549;
squeal_samples[12758]=32640;
squeal_samples[12759]=34631;
squeal_samples[12760]=36543;
squeal_samples[12761]=38362;
squeal_samples[12762]=40111;
squeal_samples[12763]=41762;
squeal_samples[12764]=43364;
squeal_samples[12765]=44868;
squeal_samples[12766]=46324;
squeal_samples[12767]=47706;
squeal_samples[12768]=49031;
squeal_samples[12769]=50296;
squeal_samples[12770]=51498;
squeal_samples[12771]=52611;
squeal_samples[12772]=49637;
squeal_samples[12773]=44401;
squeal_samples[12774]=39486;
squeal_samples[12775]=34900;
squeal_samples[12776]=30596;
squeal_samples[12777]=26579;
squeal_samples[12778]=22815;
squeal_samples[12779]=19296;
squeal_samples[12780]=15994;
squeal_samples[12781]=12920;
squeal_samples[12782]=10030;
squeal_samples[12783]=7340;
squeal_samples[12784]=7635;
squeal_samples[12785]=10720;
squeal_samples[12786]=13680;
squeal_samples[12787]=16506;
squeal_samples[12788]=19213;
squeal_samples[12789]=21802;
squeal_samples[12790]=24277;
squeal_samples[12791]=26639;
squeal_samples[12792]=28900;
squeal_samples[12793]=31064;
squeal_samples[12794]=33128;
squeal_samples[12795]=35106;
squeal_samples[12796]=36988;
squeal_samples[12797]=38789;
squeal_samples[12798]=40516;
squeal_samples[12799]=42155;
squeal_samples[12800]=43727;
squeal_samples[12801]=45229;
squeal_samples[12802]=46658;
squeal_samples[12803]=48030;
squeal_samples[12804]=49338;
squeal_samples[12805]=50589;
squeal_samples[12806]=51779;
squeal_samples[12807]=52454;
squeal_samples[12808]=48282;
squeal_samples[12809]=43122;
squeal_samples[12810]=38298;
squeal_samples[12811]=33777;
squeal_samples[12812]=29555;
squeal_samples[12813]=25598;
squeal_samples[12814]=21897;
squeal_samples[12815]=18437;
squeal_samples[12816]=15195;
squeal_samples[12817]=12162;
squeal_samples[12818]=9329;
squeal_samples[12819]=6855;
squeal_samples[12820]=8408;
squeal_samples[12821]=11459;
squeal_samples[12822]=14378;
squeal_samples[12823]=17179;
squeal_samples[12824]=19853;
squeal_samples[12825]=22417;
squeal_samples[12826]=24866;
squeal_samples[12827]=27198;
squeal_samples[12828]=29436;
squeal_samples[12829]=31573;
squeal_samples[12830]=33620;
squeal_samples[12831]=35568;
squeal_samples[12832]=37434;
squeal_samples[12833]=39215;
squeal_samples[12834]=40919;
squeal_samples[12835]=42541;
squeal_samples[12836]=44095;
squeal_samples[12837]=45574;
squeal_samples[12838]=46994;
squeal_samples[12839]=48346;
squeal_samples[12840]=49637;
squeal_samples[12841]=50881;
squeal_samples[12842]=52057;
squeal_samples[12843]=51886;
squeal_samples[12844]=46941;
squeal_samples[12845]=41875;
squeal_samples[12846]=37124;
squeal_samples[12847]=32684;
squeal_samples[12848]=28522;
squeal_samples[12849]=24641;
squeal_samples[12850]=20996;
squeal_samples[12851]=17592;
squeal_samples[12852]=14403;
squeal_samples[12853]=11420;
squeal_samples[12854]=8633;
squeal_samples[12855]=6739;
squeal_samples[12856]=9165;
squeal_samples[12857]=12188;
squeal_samples[12858]=15076;
squeal_samples[12859]=17848;
squeal_samples[12860]=20490;
squeal_samples[12861]=23027;
squeal_samples[12862]=25447;
squeal_samples[12863]=27755;
squeal_samples[12864]=29969;
squeal_samples[12865]=32079;
squeal_samples[12866]=34099;
squeal_samples[12867]=36031;
squeal_samples[12868]=37870;
squeal_samples[12869]=39634;
squeal_samples[12870]=41317;
squeal_samples[12871]=42922;
squeal_samples[12872]=44461;
squeal_samples[12873]=45923;
squeal_samples[12874]=47327;
squeal_samples[12875]=48661;
squeal_samples[12876]=49941;
squeal_samples[12877]=51162;
squeal_samples[12878]=52329;
squeal_samples[12879]=50908;
squeal_samples[12880]=45628;
squeal_samples[12881]=40642;
squeal_samples[12882]=35972;
squeal_samples[12883]=31601;
squeal_samples[12884]=27513;
squeal_samples[12885]=23688;
squeal_samples[12886]=20110;
squeal_samples[12887]=16755;
squeal_samples[12888]=13624;
squeal_samples[12889]=10693;
squeal_samples[12890]=7950;
squeal_samples[12891]=6980;
squeal_samples[12892]=9917;
squeal_samples[12893]=12906;
squeal_samples[12894]=15768;
squeal_samples[12895]=18507;
squeal_samples[12896]=21121;
squeal_samples[12897]=23627;
squeal_samples[12898]=26012;
squeal_samples[12899]=28305;
squeal_samples[12900]=30492;
squeal_samples[12901]=32580;
squeal_samples[12902]=34573;
squeal_samples[12903]=36482;
squeal_samples[12904]=38306;
squeal_samples[12905]=40050;
squeal_samples[12906]=41706;
squeal_samples[12907]=43303;
squeal_samples[12908]=44809;
squeal_samples[12909]=46266;
squeal_samples[12910]=47647;
squeal_samples[12911]=48974;
squeal_samples[12912]=50233;
squeal_samples[12913]=51444;
squeal_samples[12914]=52594;
squeal_samples[12915]=50396;
squeal_samples[12916]=45095;
squeal_samples[12917]=40147;
squeal_samples[12918]=35501;
squeal_samples[12919]=31170;
squeal_samples[12920]=27094;
squeal_samples[12921]=23306;
squeal_samples[12922]=19742;
squeal_samples[12923]=16420;
squeal_samples[12924]=13301;
squeal_samples[12925]=10394;
squeal_samples[12926]=7672;
squeal_samples[12927]=6717;
squeal_samples[12928]=9664;
squeal_samples[12929]=12663;
squeal_samples[12930]=15532;
squeal_samples[12931]=18278;
squeal_samples[12932]=20909;
squeal_samples[12933]=23419;
squeal_samples[12934]=25817;
squeal_samples[12935]=28108;
squeal_samples[12936]=30311;
squeal_samples[12937]=32402;
squeal_samples[12938]=34407;
squeal_samples[12939]=36321;
squeal_samples[12940]=38151;
squeal_samples[12941]=39897;
squeal_samples[12942]=41570;
squeal_samples[12943]=43160;
squeal_samples[12944]=44684;
squeal_samples[12945]=46142;
squeal_samples[12946]=47528;
squeal_samples[12947]=48857;
squeal_samples[12948]=50121;
squeal_samples[12949]=51334;
squeal_samples[12950]=52499;
squeal_samples[12951]=50292;
squeal_samples[12952]=45012;
squeal_samples[12953]=40049;
squeal_samples[12954]=35423;
squeal_samples[12955]=31083;
squeal_samples[12956]=27026;
squeal_samples[12957]=23231;
squeal_samples[12958]=19684;
squeal_samples[12959]=16351;
squeal_samples[12960]=13247;
squeal_samples[12961]=10338;
squeal_samples[12962]=7614;
squeal_samples[12963]=7235;
squeal_samples[12964]=10289;
squeal_samples[12965]=13263;
squeal_samples[12966]=16104;
squeal_samples[12967]=18828;
squeal_samples[12968]=21430;
squeal_samples[12969]=23917;
squeal_samples[12970]=26293;
squeal_samples[12971]=28568;
squeal_samples[12972]=30740;
squeal_samples[12973]=32817;
squeal_samples[12974]=34803;
squeal_samples[12975]=36699;
squeal_samples[12976]=38508;
squeal_samples[12977]=40244;
squeal_samples[12978]=41890;
squeal_samples[12979]=43470;
squeal_samples[12980]=44981;
squeal_samples[12981]=46423;
squeal_samples[12982]=47799;
squeal_samples[12983]=49112;
squeal_samples[12984]=50368;
squeal_samples[12985]=51570;
squeal_samples[12986]=52667;
squeal_samples[12987]=49688;
squeal_samples[12988]=44440;
squeal_samples[12989]=39521;
squeal_samples[12990]=34922;
squeal_samples[12991]=30615;
squeal_samples[12992]=26586;
squeal_samples[12993]=22821;
squeal_samples[12994]=19294;
squeal_samples[12995]=15994;
squeal_samples[12996]=12907;
squeal_samples[12997]=10019;
squeal_samples[12998]=7317;
squeal_samples[12999]=7611;
squeal_samples[13000]=10694;
squeal_samples[13001]=13650;
squeal_samples[13002]=16474;
squeal_samples[13003]=19178;
squeal_samples[13004]=21770;
squeal_samples[13005]=24236;
squeal_samples[13006]=26601;
squeal_samples[13007]=28856;
squeal_samples[13008]=31020;
squeal_samples[13009]=33083;
squeal_samples[13010]=35057;
squeal_samples[13011]=36937;
squeal_samples[13012]=38739;
squeal_samples[13013]=40463;
squeal_samples[13014]=42096;
squeal_samples[13015]=43676;
squeal_samples[13016]=45170;
squeal_samples[13017]=46601;
squeal_samples[13018]=47966;
squeal_samples[13019]=49279;
squeal_samples[13020]=50521;
squeal_samples[13021]=51719;
squeal_samples[13022]=52649;
squeal_samples[13023]=49014;
squeal_samples[13024]=43807;
squeal_samples[13025]=38925;
squeal_samples[13026]=34364;
squeal_samples[13027]=30097;
squeal_samples[13028]=26097;
squeal_samples[13029]=22364;
squeal_samples[13030]=18864;
squeal_samples[13031]=15591;
squeal_samples[13032]=12526;
squeal_samples[13033]=9663;
squeal_samples[13034]=7031;
squeal_samples[13035]=7994;
squeal_samples[13036]=11060;
squeal_samples[13037]=13998;
squeal_samples[13038]=16809;
squeal_samples[13039]=19498;
squeal_samples[13040]=22077;
squeal_samples[13041]=24532;
squeal_samples[13042]=26878;
squeal_samples[13043]=29126;
squeal_samples[13044]=31274;
squeal_samples[13045]=33325;
squeal_samples[13046]=35287;
squeal_samples[13047]=37155;
squeal_samples[13048]=38950;
squeal_samples[13049]=40656;
squeal_samples[13050]=42292;
squeal_samples[13051]=43849;
squeal_samples[13052]=45341;
squeal_samples[13053]=46765;
squeal_samples[13054]=48122;
squeal_samples[13055]=49420;
squeal_samples[13056]=50666;
squeal_samples[13057]=51851;
squeal_samples[13058]=52515;
squeal_samples[13059]=48331;
squeal_samples[13060]=43169;
squeal_samples[13061]=38327;
squeal_samples[13062]=33805;
squeal_samples[13063]=29563;
squeal_samples[13064]=25607;
squeal_samples[13065]=21898;
squeal_samples[13066]=18426;
squeal_samples[13067]=15187;
squeal_samples[13068]=12146;
squeal_samples[13069]=9308;
squeal_samples[13070]=6825;
squeal_samples[13071]=8371;
squeal_samples[13072]=11421;
squeal_samples[13073]=14343;
squeal_samples[13074]=17141;
squeal_samples[13075]=19811;
squeal_samples[13076]=22370;
squeal_samples[13077]=24818;
squeal_samples[13078]=27151;
squeal_samples[13079]=29382;
squeal_samples[13080]=31522;
squeal_samples[13081]=33559;
squeal_samples[13082]=35512;
squeal_samples[13083]=37368;
squeal_samples[13084]=39153;
squeal_samples[13085]=40848;
squeal_samples[13086]=42480;
squeal_samples[13087]=44022;
squeal_samples[13088]=45507;
squeal_samples[13089]=46924;
squeal_samples[13090]=48277;
squeal_samples[13091]=49569;
squeal_samples[13092]=50803;
squeal_samples[13093]=51979;
squeal_samples[13094]=52277;
squeal_samples[13095]=47650;
squeal_samples[13096]=42528;
squeal_samples[13097]=37733;
squeal_samples[13098]=33247;
squeal_samples[13099]=29043;
squeal_samples[13100]=25123;
squeal_samples[13101]=21435;
squeal_samples[13102]=17996;
squeal_samples[13103]=14780;
squeal_samples[13104]=11764;
squeal_samples[13105]=8950;
squeal_samples[13106]=6714;
squeal_samples[13107]=8748;
squeal_samples[13108]=11781;
squeal_samples[13109]=14689;
squeal_samples[13110]=17465;
squeal_samples[13111]=20128;
squeal_samples[13112]=22666;
squeal_samples[13113]=25106;
squeal_samples[13114]=27417;
squeal_samples[13115]=29646;
squeal_samples[13116]=31766;
squeal_samples[13117]=33798;
squeal_samples[13118]=35732;
squeal_samples[13119]=37587;
squeal_samples[13120]=39352;
squeal_samples[13121]=41047;
squeal_samples[13122]=42660;
squeal_samples[13123]=44199;
squeal_samples[13124]=45677;
squeal_samples[13125]=47084;
squeal_samples[13126]=48424;
squeal_samples[13127]=49713;
squeal_samples[13128]=50937;
squeal_samples[13129]=52110;
squeal_samples[13130]=51934;
squeal_samples[13131]=46976;
squeal_samples[13132]=41901;
squeal_samples[13133]=37138;
squeal_samples[13134]=32694;
squeal_samples[13135]=28520;
squeal_samples[13136]=24628;
squeal_samples[13137]=20985;
squeal_samples[13138]=17566;
squeal_samples[13139]=14376;
squeal_samples[13140]=11391;
squeal_samples[13141]=8598;
squeal_samples[13142]=6695;
squeal_samples[13143]=9119;
squeal_samples[13144]=12137;
squeal_samples[13145]=15027;
squeal_samples[13146]=17790;
squeal_samples[13147]=20436;
squeal_samples[13148]=22965;
squeal_samples[13149]=25381;
squeal_samples[13150]=27687;
squeal_samples[13151]=29898;
squeal_samples[13152]=32012;
squeal_samples[13153]=34028;
squeal_samples[13154]=35952;
squeal_samples[13155]=37799;
squeal_samples[13156]=39556;
squeal_samples[13157]=41240;
squeal_samples[13158]=42840;
squeal_samples[13159]=44376;
squeal_samples[13160]=45842;
squeal_samples[13161]=47238;
squeal_samples[13162]=48573;
squeal_samples[13163]=49852;
squeal_samples[13164]=51073;
squeal_samples[13165]=52241;
squeal_samples[13166]=51487;
squeal_samples[13167]=46314;
squeal_samples[13168]=41268;
squeal_samples[13169]=36558;
squeal_samples[13170]=32139;
squeal_samples[13171]=28008;
squeal_samples[13172]=24147;
squeal_samples[13173]=20528;
squeal_samples[13174]=17150;
squeal_samples[13175]=13977;
squeal_samples[13176]=11016;
squeal_samples[13177]=8245;
squeal_samples[13178]=6763;
squeal_samples[13179]=9491;
squeal_samples[13180]=12493;
squeal_samples[13181]=15365;
squeal_samples[13182]=18114;
squeal_samples[13183]=20742;
squeal_samples[13184]=23259;
squeal_samples[13185]=25661;
squeal_samples[13186]=27956;
squeal_samples[13187]=30153;
squeal_samples[13188]=32256;
squeal_samples[13189]=34260;
squeal_samples[13190]=36180;
squeal_samples[13191]=38005;
squeal_samples[13192]=39756;
squeal_samples[13193]=41425;
squeal_samples[13194]=43021;
squeal_samples[13195]=44548;
squeal_samples[13196]=46000;
squeal_samples[13197]=47400;
squeal_samples[13198]=48720;
squeal_samples[13199]=49996;
squeal_samples[13200]=51207;
squeal_samples[13201]=52368;
squeal_samples[13202]=50934;
squeal_samples[13203]=45655;
squeal_samples[13204]=40649;
squeal_samples[13205]=35976;
squeal_samples[13206]=31591;
squeal_samples[13207]=27495;
squeal_samples[13208]=23666;
squeal_samples[13209]=20080;
squeal_samples[13210]=16721;
squeal_samples[13211]=13579;
squeal_samples[13212]=10648;
squeal_samples[13213]=7894;
squeal_samples[13214]=6923;
squeal_samples[13215]=9858;
squeal_samples[13216]=12842;
squeal_samples[13217]=15699;
squeal_samples[13218]=18436;
squeal_samples[13219]=21048;
squeal_samples[13220]=23551;
squeal_samples[13221]=25939;
squeal_samples[13222]=28223;
squeal_samples[13223]=30407;
squeal_samples[13224]=32494;
squeal_samples[13225]=34494;
squeal_samples[13226]=36397;
squeal_samples[13227]=38214;
squeal_samples[13228]=39960;
squeal_samples[13229]=41613;
squeal_samples[13230]=43209;
squeal_samples[13231]=44712;
squeal_samples[13232]=46171;
squeal_samples[13233]=47549;
squeal_samples[13234]=48873;
squeal_samples[13235]=50131;
squeal_samples[13236]=51341;
squeal_samples[13237]=52494;
squeal_samples[13238]=51057;
squeal_samples[13239]=45764;
squeal_samples[13240]=40752;
squeal_samples[13241]=36067;
squeal_samples[13242]=31683;
squeal_samples[13243]=27578;
squeal_samples[13244]=23743;
squeal_samples[13245]=20151;
squeal_samples[13246]=16785;
squeal_samples[13247]=13645;
squeal_samples[13248]=10696;
squeal_samples[13249]=7949;
squeal_samples[13250]=6484;
squeal_samples[13251]=9219;
squeal_samples[13252]=12232;
squeal_samples[13253]=15114;
squeal_samples[13254]=17874;
squeal_samples[13255]=20513;
squeal_samples[13256]=23038;
squeal_samples[13257]=25451;
squeal_samples[13258]=27757;
squeal_samples[13259]=29955;
squeal_samples[13260]=32065;
squeal_samples[13261]=34077;
squeal_samples[13262]=36002;
squeal_samples[13263]=37840;
squeal_samples[13264]=39595;
squeal_samples[13265]=41272;
squeal_samples[13266]=42876;
squeal_samples[13267]=44403;
squeal_samples[13268]=45866;
squeal_samples[13269]=47262;
squeal_samples[13270]=48588;
squeal_samples[13271]=49873;
squeal_samples[13272]=51082;
squeal_samples[13273]=52256;
squeal_samples[13274]=51492;
squeal_samples[13275]=46316;
squeal_samples[13276]=41271;
squeal_samples[13277]=36552;
squeal_samples[13278]=32136;
squeal_samples[13279]=27755;
squeal_samples[13280]=23668;
squeal_samples[13281]=20083;
squeal_samples[13282]=16720;
squeal_samples[13283]=13584;
squeal_samples[13284]=10642;
squeal_samples[13285]=7897;
squeal_samples[13286]=6914;
squeal_samples[13287]=9852;
squeal_samples[13288]=12837;
squeal_samples[13289]=15692;
squeal_samples[13290]=18425;
squeal_samples[13291]=21042;
squeal_samples[13292]=23537;
squeal_samples[13293]=25929;
squeal_samples[13294]=28211;
squeal_samples[13295]=30395;
squeal_samples[13296]=32485;
squeal_samples[13297]=34474;
squeal_samples[13298]=36380;
squeal_samples[13299]=38203;
squeal_samples[13300]=39941;
squeal_samples[13301]=41601;
squeal_samples[13302]=43186;
squeal_samples[13303]=44699;
squeal_samples[13304]=46151;
squeal_samples[13305]=47533;
squeal_samples[13306]=48856;
squeal_samples[13307]=50114;
squeal_samples[13308]=51323;
squeal_samples[13309]=52473;
squeal_samples[13310]=51033;
squeal_samples[13311]=45742;
squeal_samples[13312]=40730;
squeal_samples[13313]=36049;
squeal_samples[13314]=31660;
squeal_samples[13315]=27556;
squeal_samples[13316]=23720;
squeal_samples[13317]=20128;
squeal_samples[13318]=16764;
squeal_samples[13319]=13619;
squeal_samples[13320]=10675;
squeal_samples[13321]=7925;
squeal_samples[13322]=6945;
squeal_samples[13323]=9876;
squeal_samples[13324]=12860;
squeal_samples[13325]=15717;
squeal_samples[13326]=18447;
squeal_samples[13327]=21065;
squeal_samples[13328]=23552;
squeal_samples[13329]=25945;
squeal_samples[13330]=28223;
squeal_samples[13331]=30409;
squeal_samples[13332]=32496;
squeal_samples[13333]=34489;
squeal_samples[13334]=36395;
squeal_samples[13335]=38209;
squeal_samples[13336]=39949;
squeal_samples[13337]=41609;
squeal_samples[13338]=43192;
squeal_samples[13339]=44711;
squeal_samples[13340]=46149;
squeal_samples[13341]=47539;
squeal_samples[13342]=48856;
squeal_samples[13343]=50118;
squeal_samples[13344]=51324;
squeal_samples[13345]=52477;
squeal_samples[13346]=51034;
squeal_samples[13347]=45742;
squeal_samples[13348]=40728;
squeal_samples[13349]=36050;
squeal_samples[13350]=31655;
squeal_samples[13351]=27554;
squeal_samples[13352]=23717;
squeal_samples[13353]=20125;
squeal_samples[13354]=16753;
squeal_samples[13355]=13616;
squeal_samples[13356]=10662;
squeal_samples[13357]=7921;
squeal_samples[13358]=6931;
squeal_samples[13359]=9873;
squeal_samples[13360]=12848;
squeal_samples[13361]=15711;
squeal_samples[13362]=18440;
squeal_samples[13363]=21050;
squeal_samples[13364]=23552;
squeal_samples[13365]=25930;
squeal_samples[13366]=28219;
squeal_samples[13367]=30398;
squeal_samples[13368]=32484;
squeal_samples[13369]=34480;
squeal_samples[13370]=36379;
squeal_samples[13371]=38199;
squeal_samples[13372]=39938;
squeal_samples[13373]=41597;
squeal_samples[13374]=43179;
squeal_samples[13375]=44694;
squeal_samples[13376]=46144;
squeal_samples[13377]=47524;
squeal_samples[13378]=48841;
squeal_samples[13379]=50107;
squeal_samples[13380]=51309;
squeal_samples[13381]=52468;
squeal_samples[13382]=51023;
squeal_samples[13383]=45728;
squeal_samples[13384]=40721;
squeal_samples[13385]=36031;
squeal_samples[13386]=31645;
squeal_samples[13387]=27537;
squeal_samples[13388]=23707;
squeal_samples[13389]=20108;
squeal_samples[13390]=16749;
squeal_samples[13391]=13597;
squeal_samples[13392]=10658;
squeal_samples[13393]=7904;
squeal_samples[13394]=6921;
squeal_samples[13395]=9862;
squeal_samples[13396]=12835;
squeal_samples[13397]=15698;
squeal_samples[13398]=18424;
squeal_samples[13399]=21040;
squeal_samples[13400]=23535;
squeal_samples[13401]=25918;
squeal_samples[13402]=28205;
squeal_samples[13403]=30384;
squeal_samples[13404]=32472;
squeal_samples[13405]=34464;
squeal_samples[13406]=36368;
squeal_samples[13407]=38187;
squeal_samples[13408]=39929;
squeal_samples[13409]=41579;
squeal_samples[13410]=43174;
squeal_samples[13411]=44684;
squeal_samples[13412]=46131;
squeal_samples[13413]=47509;
squeal_samples[13414]=48829;
squeal_samples[13415]=50092;
squeal_samples[13416]=51296;
squeal_samples[13417]=52454;
squeal_samples[13418]=51009;
squeal_samples[13419]=45715;
squeal_samples[13420]=40708;
squeal_samples[13421]=36016;
squeal_samples[13422]=31633;
squeal_samples[13423]=27522;
squeal_samples[13424]=23694;
squeal_samples[13425]=20094;
squeal_samples[13426]=16736;
squeal_samples[13427]=13582;
squeal_samples[13428]=10647;
squeal_samples[13429]=7888;
squeal_samples[13430]=6909;
squeal_samples[13431]=9847;
squeal_samples[13432]=12823;
squeal_samples[13433]=15682;
squeal_samples[13434]=18413;
squeal_samples[13435]=21025;
squeal_samples[13436]=23522;
squeal_samples[13437]=25905;
squeal_samples[13438]=28190;
squeal_samples[13439]=30371;
squeal_samples[13440]=32457;
squeal_samples[13441]=34453;
squeal_samples[13442]=36352;
squeal_samples[13443]=38177;
squeal_samples[13444]=39911;
squeal_samples[13445]=41574;
squeal_samples[13446]=43157;
squeal_samples[13447]=44674;
squeal_samples[13448]=46115;
squeal_samples[13449]=47497;
squeal_samples[13450]=48815;
squeal_samples[13451]=50077;
squeal_samples[13452]=51285;
squeal_samples[13453]=52438;
squeal_samples[13454]=50997;
squeal_samples[13455]=45701;
squeal_samples[13456]=40693;
squeal_samples[13457]=36005;
squeal_samples[13458]=31617;
squeal_samples[13459]=27510;
squeal_samples[13460]=23680;
squeal_samples[13461]=20080;
squeal_samples[13462]=16723;
squeal_samples[13463]=13569;
squeal_samples[13464]=10632;
squeal_samples[13465]=7876;
squeal_samples[13466]=6894;
squeal_samples[13467]=9834;
squeal_samples[13468]=12811;
squeal_samples[13469]=15666;
squeal_samples[13470]=18402;
squeal_samples[13471]=21009;
squeal_samples[13472]=23509;
squeal_samples[13473]=25893;
squeal_samples[13474]=28174;
squeal_samples[13475]=30362;
squeal_samples[13476]=32439;
squeal_samples[13477]=34442;
squeal_samples[13478]=36336;
squeal_samples[13479]=38166;
squeal_samples[13480]=39896;
squeal_samples[13481]=41563;
squeal_samples[13482]=43141;
squeal_samples[13483]=44662;
squeal_samples[13484]=46100;
squeal_samples[13485]=47485;
squeal_samples[13486]=48801;
squeal_samples[13487]=50064;
squeal_samples[13488]=51271;
squeal_samples[13489]=52425;
squeal_samples[13490]=50983;
squeal_samples[13491]=45688;
squeal_samples[13492]=40679;
squeal_samples[13493]=35992;
squeal_samples[13494]=31603;
squeal_samples[13495]=27498;
squeal_samples[13496]=23664;
squeal_samples[13497]=20068;
squeal_samples[13498]=16709;
squeal_samples[13499]=13555;
squeal_samples[13500]=10621;
squeal_samples[13501]=7858;
squeal_samples[13502]=6885;
squeal_samples[13503]=9817;
squeal_samples[13504]=12800;
squeal_samples[13505]=15652;
squeal_samples[13506]=18387;
squeal_samples[13507]=20997;
squeal_samples[13508]=23496;
squeal_samples[13509]=25878;
squeal_samples[13510]=28162;
squeal_samples[13511]=30346;
squeal_samples[13512]=32429;
squeal_samples[13513]=34426;
squeal_samples[13514]=36326;
squeal_samples[13515]=38147;
squeal_samples[13516]=39888;
squeal_samples[13517]=41544;
squeal_samples[13518]=43134;
squeal_samples[13519]=44642;
squeal_samples[13520]=46093;
squeal_samples[13521]=47467;
squeal_samples[13522]=48789;
squeal_samples[13523]=50051;
squeal_samples[13524]=51256;
squeal_samples[13525]=52413;
squeal_samples[13526]=50969;
squeal_samples[13527]=45675;
squeal_samples[13528]=40666;
squeal_samples[13529]=35977;
squeal_samples[13530]=31591;
squeal_samples[13531]=27484;
squeal_samples[13532]=23651;
squeal_samples[13533]=20055;
squeal_samples[13534]=16695;
squeal_samples[13535]=13542;
squeal_samples[13536]=10607;
squeal_samples[13537]=7846;
squeal_samples[13538]=6870;
squeal_samples[13539]=9805;
squeal_samples[13540]=12785;
squeal_samples[13541]=15639;
squeal_samples[13542]=18376;
squeal_samples[13543]=20980;
squeal_samples[13544]=23486;
squeal_samples[13545]=25860;
squeal_samples[13546]=28153;
squeal_samples[13547]=30330;
squeal_samples[13548]=32417;
squeal_samples[13549]=34412;
squeal_samples[13550]=36312;
squeal_samples[13551]=38135;
squeal_samples[13552]=39872;
squeal_samples[13553]=41535;
squeal_samples[13554]=43114;
squeal_samples[13555]=44638;
squeal_samples[13556]=46070;
squeal_samples[13557]=47460;
squeal_samples[13558]=48773;
squeal_samples[13559]=50037;
squeal_samples[13560]=51245;
squeal_samples[13561]=52399;
squeal_samples[13562]=50954;
squeal_samples[13563]=45663;
squeal_samples[13564]=40650;
squeal_samples[13565]=35967;
squeal_samples[13566]=31576;
squeal_samples[13567]=27470;
squeal_samples[13568]=23639;
squeal_samples[13569]=20039;
squeal_samples[13570]=16683;
squeal_samples[13571]=13529;
squeal_samples[13572]=10592;
squeal_samples[13573]=7835;
squeal_samples[13574]=6855;
squeal_samples[13575]=9791;
squeal_samples[13576]=12773;
squeal_samples[13577]=15625;
squeal_samples[13578]=18362;
squeal_samples[13579]=20968;
squeal_samples[13580]=23470;
squeal_samples[13581]=25850;
squeal_samples[13582]=28137;
squeal_samples[13583]=30318;
squeal_samples[13584]=32402;
squeal_samples[13585]=34399;
squeal_samples[13586]=36299;
squeal_samples[13587]=38121;
squeal_samples[13588]=39860;
squeal_samples[13589]=41519;
squeal_samples[13590]=43103;
squeal_samples[13591]=44621;
squeal_samples[13592]=46059;
squeal_samples[13593]=47446;
squeal_samples[13594]=48759;
squeal_samples[13595]=50024;
squeal_samples[13596]=51230;
squeal_samples[13597]=52383;
squeal_samples[13598]=51613;
squeal_samples[13599]=46417;
squeal_samples[13600]=41364;
squeal_samples[13601]=36627;
squeal_samples[13602]=32200;
squeal_samples[13603]=28055;
squeal_samples[13604]=24176;
squeal_samples[13605]=20552;
squeal_samples[13606]=17149;
squeal_samples[13607]=13974;
squeal_samples[13608]=11000;
squeal_samples[13609]=8225;
squeal_samples[13610]=6731;
squeal_samples[13611]=9456;
squeal_samples[13612]=12445;
squeal_samples[13613]=15315;
squeal_samples[13614]=18059;
squeal_samples[13615]=20685;
squeal_samples[13616]=23195;
squeal_samples[13617]=25594;
squeal_samples[13618]=27882;
squeal_samples[13619]=30080;
squeal_samples[13620]=32173;
squeal_samples[13621]=34184;
squeal_samples[13622]=36086;
squeal_samples[13623]=37921;
squeal_samples[13624]=39660;
squeal_samples[13625]=41332;
squeal_samples[13626]=42923;
squeal_samples[13627]=44447;
squeal_samples[13628]=45898;
squeal_samples[13629]=47286;
squeal_samples[13630]=48615;
squeal_samples[13631]=49876;
squeal_samples[13632]=51094;
squeal_samples[13633]=52248;
squeal_samples[13634]=52058;
squeal_samples[13635]=47081;
squeal_samples[13636]=41987;
squeal_samples[13637]=37206;
squeal_samples[13638]=32740;
squeal_samples[13639]=28557;
squeal_samples[13640]=24654;
squeal_samples[13641]=20986;
squeal_samples[13642]=17561;
squeal_samples[13643]=14357;
squeal_samples[13644]=11356;
squeal_samples[13645]=8560;
squeal_samples[13646]=6643;
squeal_samples[13647]=9064;
squeal_samples[13648]=12074;
squeal_samples[13649]=14963;
squeal_samples[13650]=17715;
squeal_samples[13651]=20361;
squeal_samples[13652]=22880;
squeal_samples[13653]=25298;
squeal_samples[13654]=27601;
squeal_samples[13655]=29801;
squeal_samples[13656]=31911;
squeal_samples[13657]=33919;
squeal_samples[13658]=35851;
squeal_samples[13659]=37681;
squeal_samples[13660]=39443;
squeal_samples[13661]=41118;
squeal_samples[13662]=42718;
squeal_samples[13663]=44251;
squeal_samples[13664]=45709;
squeal_samples[13665]=47107;
squeal_samples[13666]=48441;
squeal_samples[13667]=49714;
squeal_samples[13668]=50930;
squeal_samples[13669]=52098;
squeal_samples[13670]=52376;
squeal_samples[13671]=47736;
squeal_samples[13672]=42589;
squeal_samples[13673]=37777;
squeal_samples[13674]=33274;
squeal_samples[13675]=29055;
squeal_samples[13676]=25111;
squeal_samples[13677]=21421;
squeal_samples[13678]=17964;
squeal_samples[13679]=14736;
squeal_samples[13680]=11712;
squeal_samples[13681]=8883;
squeal_samples[13682]=6642;
squeal_samples[13683]=8663;
squeal_samples[13684]=11695;
squeal_samples[13685]=14591;
squeal_samples[13686]=17371;
squeal_samples[13687]=20022;
squeal_samples[13688]=22562;
squeal_samples[13689]=24984;
squeal_samples[13690]=27306;
squeal_samples[13691]=29516;
squeal_samples[13692]=31643;
squeal_samples[13693]=33662;
squeal_samples[13694]=35603;
squeal_samples[13695]=37448;
squeal_samples[13696]=39210;
squeal_samples[13697]=40900;
squeal_samples[13698]=42510;
squeal_samples[13699]=44051;
squeal_samples[13700]=45520;
squeal_samples[13701]=46922;
squeal_samples[13702]=48268;
squeal_samples[13703]=49546;
squeal_samples[13704]=50772;
squeal_samples[13705]=51941;
squeal_samples[13706]=52593;
squeal_samples[13707]=48390;
squeal_samples[13708]=43201;
squeal_samples[13709]=38349;
squeal_samples[13710]=33806;
squeal_samples[13711]=29550;
squeal_samples[13712]=25579;
squeal_samples[13713]=21855;
squeal_samples[13714]=18377;
squeal_samples[13715]=15111;
squeal_samples[13716]=12066;
squeal_samples[13717]=9215;
squeal_samples[13718]=6729;
squeal_samples[13719]=8262;
squeal_samples[13720]=11312;
squeal_samples[13721]=14226;
squeal_samples[13722]=17014;
squeal_samples[13723]=19686;
squeal_samples[13724]=22237;
squeal_samples[13725]=24678;
squeal_samples[13726]=27012;
squeal_samples[13727]=29229;
squeal_samples[13728]=31371;
squeal_samples[13729]=33400;
squeal_samples[13730]=35351;
squeal_samples[13731]=37205;
squeal_samples[13732]=38987;
squeal_samples[13733]=40679;
squeal_samples[13734]=42302;
squeal_samples[13735]=43850;
squeal_samples[13736]=45324;
squeal_samples[13737]=46738;
squeal_samples[13738]=48090;
squeal_samples[13739]=49376;
squeal_samples[13740]=50607;
squeal_samples[13741]=51786;
squeal_samples[13742]=52704;
squeal_samples[13743]=49045;
squeal_samples[13744]=43819;
squeal_samples[13745]=38923;
squeal_samples[13746]=34344;
squeal_samples[13747]=30063;
squeal_samples[13748]=26043;
squeal_samples[13749]=22298;
squeal_samples[13750]=18779;
squeal_samples[13751]=15496;
squeal_samples[13752]=12421;
squeal_samples[13753]=9546;
squeal_samples[13754]=6903;
squeal_samples[13755]=7862;
squeal_samples[13756]=10921;
squeal_samples[13757]=13855;
squeal_samples[13758]=16660;
squeal_samples[13759]=19345;
squeal_samples[13760]=21909;
squeal_samples[13761]=24369;
squeal_samples[13762]=26706;
squeal_samples[13763]=28951;
squeal_samples[13764]=31093;
squeal_samples[13765]=33138;
squeal_samples[13766]=35099;
squeal_samples[13767]=36964;
squeal_samples[13768]=38758;
squeal_samples[13769]=40458;
squeal_samples[13770]=42090;
squeal_samples[13771]=43644;
squeal_samples[13772]=45134;
squeal_samples[13773]=46551;
squeal_samples[13774]=47907;
squeal_samples[13775]=49208;
squeal_samples[13776]=50445;
squeal_samples[13777]=51626;
squeal_samples[13778]=52707;
squeal_samples[13779]=49711;
squeal_samples[13780]=44444;
squeal_samples[13781]=39504;
squeal_samples[13782]=34890;
squeal_samples[13783]=30559;
squeal_samples[13784]=26520;
squeal_samples[13785]=22736;
squeal_samples[13786]=19198;
squeal_samples[13787]=15884;
squeal_samples[13788]=12783;
squeal_samples[13789]=9880;
squeal_samples[13790]=7174;
squeal_samples[13791]=7456;
squeal_samples[13792]=10533;
squeal_samples[13793]=13485;
squeal_samples[13794]=16303;
squeal_samples[13795]=19001;
squeal_samples[13796]=21583;
squeal_samples[13797]=24048;
squeal_samples[13798]=26409;
squeal_samples[13799]=28659;
squeal_samples[13800]=30820;
squeal_samples[13801]=32876;
squeal_samples[13802]=34846;
squeal_samples[13803]=36725;
squeal_samples[13804]=38519;
squeal_samples[13805]=40237;
squeal_samples[13806]=41873;
squeal_samples[13807]=43444;
squeal_samples[13808]=44935;
squeal_samples[13809]=46364;
squeal_samples[13810]=47731;
squeal_samples[13811]=49037;
squeal_samples[13812]=50280;
squeal_samples[13813]=51472;
squeal_samples[13814]=52611;
squeal_samples[13815]=50384;
squeal_samples[13816]=45069;
squeal_samples[13817]=40092;
squeal_samples[13818]=35438;
squeal_samples[13819]=31076;
squeal_samples[13820]=26999;
squeal_samples[13821]=23186;
squeal_samples[13822]=19612;
squeal_samples[13823]=16274;
squeal_samples[13824]=13144;
squeal_samples[13825]=10222;
squeal_samples[13826]=7486;
squeal_samples[13827]=7094;
squeal_samples[13828]=10147;
squeal_samples[13829]=13105;
squeal_samples[13830]=15945;
squeal_samples[13831]=18655;
squeal_samples[13832]=21255;
squeal_samples[13833]=23733;
squeal_samples[13834]=26107;
squeal_samples[13835]=28374;
squeal_samples[13836]=30541;
squeal_samples[13837]=32614;
squeal_samples[13838]=34588;
squeal_samples[13839]=36486;
squeal_samples[13840]=38287;
squeal_samples[13841]=40019;
squeal_samples[13842]=41658;
squeal_samples[13843]=43236;
squeal_samples[13844]=44743;
squeal_samples[13845]=46177;
squeal_samples[13846]=47550;
squeal_samples[13847]=48861;
squeal_samples[13848]=50114;
squeal_samples[13849]=51313;
squeal_samples[13850]=52455;
squeal_samples[13851]=51008;
squeal_samples[13852]=45703;
squeal_samples[13853]=40681;
squeal_samples[13854]=35991;
squeal_samples[13855]=31589;
squeal_samples[13856]=27480;
squeal_samples[13857]=23636;
squeal_samples[13858]=20032;
squeal_samples[13859]=16669;
squeal_samples[13860]=13511;
squeal_samples[13861]=10568;
squeal_samples[13862]=7804;
squeal_samples[13863]=6822;
squeal_samples[13864]=9750;
squeal_samples[13865]=12732;
squeal_samples[13866]=15581;
squeal_samples[13867]=18314;
squeal_samples[13868]=20924;
squeal_samples[13869]=23418;
squeal_samples[13870]=25800;
squeal_samples[13871]=28079;
squeal_samples[13872]=30264;
squeal_samples[13873]=32342;
squeal_samples[13874]=34341;
squeal_samples[13875]=36234;
squeal_samples[13876]=38056;
squeal_samples[13877]=39791;
squeal_samples[13878]=41448;
squeal_samples[13879]=43029;
squeal_samples[13880]=44549;
squeal_samples[13881]=45987;
squeal_samples[13882]=47371;
squeal_samples[13883]=48688;
squeal_samples[13884]=49951;
squeal_samples[13885]=51152;
squeal_samples[13886]=52301;
squeal_samples[13887]=51532;
squeal_samples[13888]=46337;
squeal_samples[13889]=41276;
squeal_samples[13890]=36548;
squeal_samples[13891]=32115;
squeal_samples[13892]=27965;
squeal_samples[13893]=24090;
squeal_samples[13894]=20455;
squeal_samples[13895]=17060;
squeal_samples[13896]=13888;
squeal_samples[13897]=10903;
squeal_samples[13898]=8133;
squeal_samples[13899]=6637;
squeal_samples[13900]=9358;
squeal_samples[13901]=12355;
squeal_samples[13902]=15219;
squeal_samples[13903]=17965;
squeal_samples[13904]=20592;
squeal_samples[13905]=23099;
squeal_samples[13906]=25495;
squeal_samples[13907]=27789;
squeal_samples[13908]=29983;
squeal_samples[13909]=32077;
squeal_samples[13910]=34080;
squeal_samples[13911]=35991;
squeal_samples[13912]=37818;
squeal_samples[13913]=39568;
squeal_samples[13914]=41231;
squeal_samples[13915]=42824;
squeal_samples[13916]=44343;
squeal_samples[13917]=45796;
squeal_samples[13918]=47190;
squeal_samples[13919]=48511;
squeal_samples[13920]=49781;
squeal_samples[13921]=50989;
squeal_samples[13922]=52149;
squeal_samples[13923]=52418;
squeal_samples[13924]=47771;
squeal_samples[13925]=42616;
squeal_samples[13926]=37798;
squeal_samples[13927]=33288;
squeal_samples[13928]=29059;
squeal_samples[13929]=25112;
squeal_samples[13930]=21417;
squeal_samples[13931]=17952;
squeal_samples[13932]=14722;
squeal_samples[13933]=11690;
squeal_samples[13934]=8858;
squeal_samples[13935]=6607;
squeal_samples[13936]=8635;
squeal_samples[13937]=11659;
squeal_samples[13938]=14557;
squeal_samples[13939]=17327;
squeal_samples[13940]=19980;
squeal_samples[13941]=22518;
squeal_samples[13942]=24944;
squeal_samples[13943]=27254;
squeal_samples[13944]=29472;
squeal_samples[13945]=31585;
squeal_samples[13946]=33613;
squeal_samples[13947]=35542;
squeal_samples[13948]=37389;
squeal_samples[13949]=39152;
squeal_samples[13950]=40838;
squeal_samples[13951]=42454;
squeal_samples[13952]=43986;
squeal_samples[13953]=45454;
squeal_samples[13954]=46861;
squeal_samples[13955]=48199;
squeal_samples[13956]=49479;
squeal_samples[13957]=50701;
squeal_samples[13958]=51871;
squeal_samples[13959]=52783;
squeal_samples[13960]=49119;
squeal_samples[13961]=43881;
squeal_samples[13962]=38976;
squeal_samples[13963]=34385;
squeal_samples[13964]=30091;
squeal_samples[13965]=26072;
squeal_samples[13966]=22318;
squeal_samples[13967]=18802;
squeal_samples[13968]=15503;
squeal_samples[13969]=12424;
squeal_samples[13970]=9544;
squeal_samples[13971]=6896;
squeal_samples[13972]=7853;
squeal_samples[13973]=10908;
squeal_samples[13974]=13838;
squeal_samples[13975]=16639;
squeal_samples[13976]=19323;
squeal_samples[13977]=21884;
squeal_samples[13978]=24340;
squeal_samples[13979]=26677;
squeal_samples[13980]=28921;
squeal_samples[13981]=31058;
squeal_samples[13982]=33104;
squeal_samples[13983]=35064;
squeal_samples[13984]=36929;
squeal_samples[13985]=38711;
squeal_samples[13986]=40419;
squeal_samples[13987]=42049;
squeal_samples[13988]=43600;
squeal_samples[13989]=45087;
squeal_samples[13990]=46505;
squeal_samples[13991]=47862;
squeal_samples[13992]=49156;
squeal_samples[13993]=50393;
squeal_samples[13994]=51577;
squeal_samples[13995]=52700;
squeal_samples[13996]=50475;
squeal_samples[13997]=45142;
squeal_samples[13998]=40165;
squeal_samples[13999]=35496;
squeal_samples[14000]=31131;
squeal_samples[14001]=27042;
squeal_samples[14002]=23223;
squeal_samples[14003]=19648;
squeal_samples[14004]=16293;
squeal_samples[14005]=13166;
squeal_samples[14006]=10239;
squeal_samples[14007]=7495;
squeal_samples[14008]=7104;
squeal_samples[14009]=10142;
squeal_samples[14010]=13109;
squeal_samples[14011]=15941;
squeal_samples[14012]=18655;
squeal_samples[14013]=21240;
squeal_samples[14014]=23725;
squeal_samples[14015]=26088;
squeal_samples[14016]=28361;
squeal_samples[14017]=30524;
squeal_samples[14018]=32591;
squeal_samples[14019]=34569;
squeal_samples[14020]=36454;
squeal_samples[14021]=38266;
squeal_samples[14022]=39981;
squeal_samples[14023]=41635;
squeal_samples[14024]=43207;
squeal_samples[14025]=44710;
squeal_samples[14026]=46146;
squeal_samples[14027]=47511;
squeal_samples[14028]=48823;
squeal_samples[14029]=50076;
squeal_samples[14030]=51275;
squeal_samples[14031]=52415;
squeal_samples[14032]=51643;
squeal_samples[14033]=46425;
squeal_samples[14034]=41370;
squeal_samples[14035]=36619;
squeal_samples[14036]=32181;
squeal_samples[14037]=28031;
squeal_samples[14038]=24142;
squeal_samples[14039]=20508;
squeal_samples[14040]=17104;
squeal_samples[14041]=13910;
squeal_samples[14042]=10941;
squeal_samples[14043]=8149;
squeal_samples[14044]=6661;
squeal_samples[14045]=9371;
squeal_samples[14046]=12366;
squeal_samples[14047]=15229;
squeal_samples[14048]=17972;
squeal_samples[14049]=20593;
squeal_samples[14050]=23105;
squeal_samples[14051]=25494;
squeal_samples[14052]=27790;
squeal_samples[14053]=29975;
squeal_samples[14054]=32074;
squeal_samples[14055]=34067;
squeal_samples[14056]=35986;
squeal_samples[14057]=37803;
squeal_samples[14058]=39548;
squeal_samples[14059]=41214;
squeal_samples[14060]=42807;
squeal_samples[14061]=44333;
squeal_samples[14062]=45774;
squeal_samples[14063]=47167;
squeal_samples[14064]=48486;
squeal_samples[14065]=49755;
squeal_samples[14066]=50967;
squeal_samples[14067]=52122;
squeal_samples[14068]=52389;
squeal_samples[14069]=47742;
squeal_samples[14070]=42584;
squeal_samples[14071]=37766;
squeal_samples[14072]=33248;
squeal_samples[14073]=29027;
squeal_samples[14074]=25076;
squeal_samples[14075]=21381;
squeal_samples[14076]=17918;
squeal_samples[14077]=14680;
squeal_samples[14078]=11649;
squeal_samples[14079]=8824;
squeal_samples[14080]=6566;
squeal_samples[14081]=8593;
squeal_samples[14082]=11615;
squeal_samples[14083]=14514;
squeal_samples[14084]=17287;
squeal_samples[14085]=19934;
squeal_samples[14086]=22472;
squeal_samples[14087]=24896;
squeal_samples[14088]=27212;
squeal_samples[14089]=29421;
squeal_samples[14090]=31544;
squeal_samples[14091]=33561;
squeal_samples[14092]=35500;
squeal_samples[14093]=37341;
squeal_samples[14094]=39111;
squeal_samples[14095]=40795;
squeal_samples[14096]=42404;
squeal_samples[14097]=43942;
squeal_samples[14098]=45408;
squeal_samples[14099]=46812;
squeal_samples[14100]=48151;
squeal_samples[14101]=49432;
squeal_samples[14102]=50654;
squeal_samples[14103]=51826;
squeal_samples[14104]=52730;
squeal_samples[14105]=49069;
squeal_samples[14106]=43829;
squeal_samples[14107]=38930;
squeal_samples[14108]=34339;
squeal_samples[14109]=30045;
squeal_samples[14110]=26024;
squeal_samples[14111]=22271;
squeal_samples[14112]=18745;
squeal_samples[14113]=15463;
squeal_samples[14114]=12373;
squeal_samples[14115]=9501;
squeal_samples[14116]=6843;
squeal_samples[14117]=7802;
squeal_samples[14118]=10862;
squeal_samples[14119]=13787;
squeal_samples[14120]=16586;
squeal_samples[14121]=19274;
squeal_samples[14122]=21836;
squeal_samples[14123]=24290;
squeal_samples[14124]=26625;
squeal_samples[14125]=28869;
squeal_samples[14126]=31013;
squeal_samples[14127]=33057;
squeal_samples[14128]=35013;
squeal_samples[14129]=36879;
squeal_samples[14130]=38664;
squeal_samples[14131]=40368;
squeal_samples[14132]=41997;
squeal_samples[14133]=43548;
squeal_samples[14134]=45038;
squeal_samples[14135]=46452;
squeal_samples[14136]=47811;
squeal_samples[14137]=49104;
squeal_samples[14138]=50342;
squeal_samples[14139]=51526;
squeal_samples[14140]=52655;
squeal_samples[14141]=50422;
squeal_samples[14142]=45091;
squeal_samples[14143]=40114;
squeal_samples[14144]=35445;
squeal_samples[14145]=31079;
squeal_samples[14146]=26991;
squeal_samples[14147]=23172;
squeal_samples[14148]=19595;
squeal_samples[14149]=16244;
squeal_samples[14150]=13114;
squeal_samples[14151]=10186;
squeal_samples[14152]=7447;
squeal_samples[14153]=7047;
squeal_samples[14154]=10098;
squeal_samples[14155]=13052;
squeal_samples[14156]=15895;
squeal_samples[14157]=18597;
squeal_samples[14158]=21195;
squeal_samples[14159]=23669;
squeal_samples[14160]=26041;
squeal_samples[14161]=28307;
squeal_samples[14162]=30472;
squeal_samples[14163]=32542;
squeal_samples[14164]=34516;
squeal_samples[14165]=36404;
squeal_samples[14166]=38214;
squeal_samples[14167]=39934;
squeal_samples[14168]=41587;
squeal_samples[14169]=43151;
squeal_samples[14170]=44665;
squeal_samples[14171]=46088;
squeal_samples[14172]=47466;
squeal_samples[14173]=48766;
squeal_samples[14174]=50031;
squeal_samples[14175]=51217;
squeal_samples[14176]=52372;
squeal_samples[14177]=51582;
squeal_samples[14178]=46383;
squeal_samples[14179]=41313;
squeal_samples[14180]=36570;
squeal_samples[14181]=32130;
squeal_samples[14182]=27978;
squeal_samples[14183]=24093;
squeal_samples[14184]=20457;
squeal_samples[14185]=17050;
squeal_samples[14186]=13862;
squeal_samples[14187]=10887;
squeal_samples[14188]=8100;
squeal_samples[14189]=6609;
squeal_samples[14190]=9320;
squeal_samples[14191]=12314;
squeal_samples[14192]=15179;
squeal_samples[14193]=17919;
squeal_samples[14194]=20545;
squeal_samples[14195]=23050;
squeal_samples[14196]=25446;
squeal_samples[14197]=27735;
squeal_samples[14198]=29930;
squeal_samples[14199]=32016;
squeal_samples[14200]=34022;
squeal_samples[14201]=35930;
squeal_samples[14202]=37755;
squeal_samples[14203]=39496;
squeal_samples[14204]=41161;
squeal_samples[14205]=42760;
squeal_samples[14206]=44276;
squeal_samples[14207]=45729;
squeal_samples[14208]=47112;
squeal_samples[14209]=48435;
squeal_samples[14210]=49706;
squeal_samples[14211]=50914;
squeal_samples[14212]=52070;
squeal_samples[14213]=52342;
squeal_samples[14214]=47686;
squeal_samples[14215]=42536;
squeal_samples[14216]=37712;
squeal_samples[14217]=33200;
squeal_samples[14218]=28974;
squeal_samples[14219]=25027;
squeal_samples[14220]=21326;
squeal_samples[14221]=17871;
squeal_samples[14222]=14625;
squeal_samples[14223]=11602;
squeal_samples[14224]=8769;
squeal_samples[14225]=6517;
squeal_samples[14226]=8542;
squeal_samples[14227]=11562;
squeal_samples[14228]=14466;
squeal_samples[14229]=17232;
squeal_samples[14230]=19887;
squeal_samples[14231]=22418;
squeal_samples[14232]=24845;
squeal_samples[14233]=27162;
squeal_samples[14234]=29369;
squeal_samples[14235]=31492;
squeal_samples[14236]=33514;
squeal_samples[14237]=35443;
squeal_samples[14238]=37295;
squeal_samples[14239]=39057;
squeal_samples[14240]=40743;
squeal_samples[14241]=42356;
squeal_samples[14242]=43888;
squeal_samples[14243]=45358;
squeal_samples[14244]=46761;
squeal_samples[14245]=48099;
squeal_samples[14246]=49380;
squeal_samples[14247]=50605;
squeal_samples[14248]=51771;
squeal_samples[14249]=52838;
squeal_samples[14250]=49827;
squeal_samples[14251]=44537;
squeal_samples[14252]=39587;
squeal_samples[14253]=34950;
squeal_samples[14254]=30611;
squeal_samples[14255]=26558;
squeal_samples[14256]=22757;
squeal_samples[14257]=19210;
squeal_samples[14258]=15879;
squeal_samples[14259]=12772;
squeal_samples[14260]=9860;
squeal_samples[14261]=7141;
squeal_samples[14262]=7419;
squeal_samples[14263]=10490;
squeal_samples[14264]=13431;
squeal_samples[14265]=16248;
squeal_samples[14266]=18944;
squeal_samples[14267]=21516;
squeal_samples[14268]=23981;
squeal_samples[14269]=26333;
squeal_samples[14270]=28582;
squeal_samples[14271]=30735;
squeal_samples[14272]=32788;
squeal_samples[14273]=34757;
squeal_samples[14274]=36630;
squeal_samples[14275]=38426;
squeal_samples[14276]=40136;
squeal_samples[14277]=41773;
squeal_samples[14278]=43334;
squeal_samples[14279]=44827;
squeal_samples[14280]=46257;
squeal_samples[14281]=47616;
squeal_samples[14282]=48920;
squeal_samples[14283]=50157;
squeal_samples[14284]=51351;
squeal_samples[14285]=52482;
squeal_samples[14286]=51697;
squeal_samples[14287]=46480;
squeal_samples[14288]=41410;
squeal_samples[14289]=36653;
squeal_samples[14290]=32207;
squeal_samples[14291]=28047;
squeal_samples[14292]=24153;
squeal_samples[14293]=20511;
squeal_samples[14294]=17098;
squeal_samples[14295]=13911;
squeal_samples[14296]=10929;
squeal_samples[14297]=8134;
squeal_samples[14298]=6635;
squeal_samples[14299]=9345;
squeal_samples[14300]=12338;
squeal_samples[14301]=15198;
squeal_samples[14302]=17943;
squeal_samples[14303]=20559;
squeal_samples[14304]=23067;
squeal_samples[14305]=25456;
squeal_samples[14306]=27745;
squeal_samples[14307]=29936;
squeal_samples[14308]=32020;
squeal_samples[14309]=34023;
squeal_samples[14310]=35929;
squeal_samples[14311]=37753;
squeal_samples[14312]=39498;
squeal_samples[14313]=41159;
squeal_samples[14314]=42755;
squeal_samples[14315]=44266;
squeal_samples[14316]=45720;
squeal_samples[14317]=47108;
squeal_samples[14318]=48423;
squeal_samples[14319]=49695;
squeal_samples[14320]=50897;
squeal_samples[14321]=52055;
squeal_samples[14322]=52685;
squeal_samples[14323]=48471;
squeal_samples[14324]=43261;
squeal_samples[14325]=38394;
squeal_samples[14326]=33827;
squeal_samples[14327]=29566;
squeal_samples[14328]=25570;
squeal_samples[14329]=21836;
squeal_samples[14330]=18342;
squeal_samples[14331]=15073;
squeal_samples[14332]=12010;
squeal_samples[14333]=9154;
squeal_samples[14334]=6648;
squeal_samples[14335]=8186;
squeal_samples[14336]=11218;
squeal_samples[14337]=14135;
squeal_samples[14338]=16912;
squeal_samples[14339]=19580;
squeal_samples[14340]=22127;
squeal_samples[14341]=24562;
squeal_samples[14342]=26889;
squeal_samples[14343]=29111;
squeal_samples[14344]=31240;
squeal_samples[14345]=33270;
squeal_samples[14346]=35211;
squeal_samples[14347]=37069;
squeal_samples[14348]=38842;
squeal_samples[14349]=40537;
squeal_samples[14350]=42153;
squeal_samples[14351]=43695;
squeal_samples[14352]=45171;
squeal_samples[14353]=46583;
squeal_samples[14354]=47924;
squeal_samples[14355]=49212;
squeal_samples[14356]=50441;
squeal_samples[14357]=51614;
squeal_samples[14358]=52740;
squeal_samples[14359]=50494;
squeal_samples[14360]=45164;
squeal_samples[14361]=40166;
squeal_samples[14362]=35493;
squeal_samples[14363]=31118;
squeal_samples[14364]=27022;
squeal_samples[14365]=23200;
squeal_samples[14366]=19616;
squeal_samples[14367]=16257;
squeal_samples[14368]=13123;
squeal_samples[14369]=10182;
squeal_samples[14370]=7444;
squeal_samples[14371]=7041;
squeal_samples[14372]=10083;
squeal_samples[14373]=13046;
squeal_samples[14374]=15873;
squeal_samples[14375]=18585;
squeal_samples[14376]=21175;
squeal_samples[14377]=23648;
squeal_samples[14378]=26014;
squeal_samples[14379]=28278;
squeal_samples[14380]=30441;
squeal_samples[14381]=32507;
squeal_samples[14382]=34484;
squeal_samples[14383]=36371;
squeal_samples[14384]=38176;
squeal_samples[14385]=39890;
squeal_samples[14386]=41542;
squeal_samples[14387]=43109;
squeal_samples[14388]=44613;
squeal_samples[14389]=46048;
squeal_samples[14390]=47418;
squeal_samples[14391]=48726;
squeal_samples[14392]=49977;
squeal_samples[14393]=51167;
squeal_samples[14394]=52311;
squeal_samples[14395]=52097;
squeal_samples[14396]=47107;
squeal_samples[14397]=41989;
squeal_samples[14398]=37198;
squeal_samples[14399]=32712;
squeal_samples[14400]=28513;
squeal_samples[14401]=24595;
squeal_samples[14402]=20915;
squeal_samples[14403]=17482;
squeal_samples[14404]=14257;
squeal_samples[14405]=11254;
squeal_samples[14406]=8442;
squeal_samples[14407]=6516;
squeal_samples[14408]=8931;
squeal_samples[14409]=11934;
squeal_samples[14410]=14812;
squeal_samples[14411]=17570;
squeal_samples[14412]=20198;
squeal_samples[14413]=22722;
squeal_samples[14414]=25129;
squeal_samples[14415]=27427;
squeal_samples[14416]=29629;
squeal_samples[14417]=31730;
squeal_samples[14418]=33738;
squeal_samples[14419]=35661;
squeal_samples[14420]=37491;
squeal_samples[14421]=39249;
squeal_samples[14422]=40915;
squeal_samples[14423]=42521;
squeal_samples[14424]=44043;
squeal_samples[14425]=45506;
squeal_samples[14426]=46898;
squeal_samples[14427]=48233;
squeal_samples[14428]=49499;
squeal_samples[14429]=50717;
squeal_samples[14430]=51876;
squeal_samples[14431]=52782;
squeal_samples[14432]=49104;
squeal_samples[14433]=43857;
squeal_samples[14434]=38945;
squeal_samples[14435]=34345;
squeal_samples[14436]=30043;
squeal_samples[14437]=26021;
squeal_samples[14438]=22256;
squeal_samples[14439]=18726;
squeal_samples[14440]=15433;
squeal_samples[14441]=12341;
squeal_samples[14442]=9463;
squeal_samples[14443]=6804;
squeal_samples[14444]=7759;
squeal_samples[14445]=10812;
squeal_samples[14446]=13738;
squeal_samples[14447]=16538;
squeal_samples[14448]=19216;
squeal_samples[14449]=21781;
squeal_samples[14450]=24224;
squeal_samples[14451]=26566;
squeal_samples[14452]=28798;
squeal_samples[14453]=30947;
squeal_samples[14454]=32981;
squeal_samples[14455]=34943;
squeal_samples[14456]=36795;
squeal_samples[14457]=38594;
squeal_samples[14458]=40283;
squeal_samples[14459]=41916;
squeal_samples[14460]=43469;
squeal_samples[14461]=44950;
squeal_samples[14462]=46377;
squeal_samples[14463]=47717;
squeal_samples[14464]=49024;
squeal_samples[14465]=50249;
squeal_samples[14466]=51441;
squeal_samples[14467]=52561;
squeal_samples[14468]=51101;
squeal_samples[14469]=45771;
squeal_samples[14470]=40737;
squeal_samples[14471]=36021;
squeal_samples[14472]=31611;
squeal_samples[14473]=27485;
squeal_samples[14474]=23623;
squeal_samples[14475]=20012;
squeal_samples[14476]=16630;
squeal_samples[14477]=13461;
squeal_samples[14478]=10507;
squeal_samples[14479]=7741;
squeal_samples[14480]=6743;
squeal_samples[14481]=9671;
squeal_samples[14482]=12642;
squeal_samples[14483]=15491;
squeal_samples[14484]=18208;
squeal_samples[14485]=20819;
squeal_samples[14486]=23306;
squeal_samples[14487]=25686;
squeal_samples[14488]=27962;
squeal_samples[14489]=30135;
squeal_samples[14490]=32216;
squeal_samples[14491]=34201;
squeal_samples[14492]=36100;
squeal_samples[14493]=37915;
squeal_samples[14494]=39643;
squeal_samples[14495]=41302;
squeal_samples[14496]=42882;
squeal_samples[14497]=44396;
squeal_samples[14498]=45830;
squeal_samples[14499]=47214;
squeal_samples[14500]=48524;
squeal_samples[14501]=49783;
squeal_samples[14502]=50981;
squeal_samples[14503]=52133;
squeal_samples[14504]=52396;
squeal_samples[14505]=47732;
squeal_samples[14506]=42572;
squeal_samples[14507]=37740;
squeal_samples[14508]=33219;
squeal_samples[14509]=28985;
squeal_samples[14510]=25035;
squeal_samples[14511]=21324;
squeal_samples[14512]=17861;
squeal_samples[14513]=14611;
squeal_samples[14514]=11582;
squeal_samples[14515]=8743;
squeal_samples[14516]=6488;
squeal_samples[14517]=8506;
squeal_samples[14518]=11525;
squeal_samples[14519]=14425;
squeal_samples[14520]=17191;
squeal_samples[14521]=19845;
squeal_samples[14522]=22372;
squeal_samples[14523]=24799;
squeal_samples[14524]=27107;
squeal_samples[14525]=29320;
squeal_samples[14526]=31439;
squeal_samples[14527]=33454;
squeal_samples[14528]=35390;
squeal_samples[14529]=37232;
squeal_samples[14530]=38993;
squeal_samples[14531]=40678;
squeal_samples[14532]=42288;
squeal_samples[14533]=43819;
squeal_samples[14534]=45291;
squeal_samples[14535]=46687;
squeal_samples[14536]=48030;
squeal_samples[14537]=49306;
squeal_samples[14538]=50531;
squeal_samples[14539]=51693;
squeal_samples[14540]=52765;
squeal_samples[14541]=49746;
squeal_samples[14542]=44454;
squeal_samples[14543]=39505;
squeal_samples[14544]=34867;
squeal_samples[14545]=30528;
squeal_samples[14546]=26470;
squeal_samples[14547]=22676;
squeal_samples[14548]=19117;
squeal_samples[14549]=15796;
squeal_samples[14550]=12681;
squeal_samples[14551]=9772;
squeal_samples[14552]=7048;
squeal_samples[14553]=7331;
squeal_samples[14554]=10400;
squeal_samples[14555]=13340;
squeal_samples[14556]=16155;
squeal_samples[14557]=18847;
squeal_samples[14558]=21426;
squeal_samples[14559]=23892;
squeal_samples[14560]=26242;
squeal_samples[14561]=28487;
squeal_samples[14562]=30646;
squeal_samples[14563]=32692;
squeal_samples[14564]=34661;
squeal_samples[14565]=36537;
squeal_samples[14566]=38327;
squeal_samples[14567]=40044;
squeal_samples[14568]=41675;
squeal_samples[14569]=43240;
squeal_samples[14570]=44733;
squeal_samples[14571]=46159;
squeal_samples[14572]=47524;
squeal_samples[14573]=48820;
squeal_samples[14574]=50067;
squeal_samples[14575]=51249;
squeal_samples[14576]=52393;
squeal_samples[14577]=52166;
squeal_samples[14578]=47172;
squeal_samples[14579]=42039;
squeal_samples[14580]=37243;
squeal_samples[14581]=32754;
squeal_samples[14582]=28547;
squeal_samples[14583]=24620;
squeal_samples[14584]=20932;
squeal_samples[14585]=17497;
squeal_samples[14586]=14268;
squeal_samples[14587]=11260;
squeal_samples[14588]=8435;
squeal_samples[14589]=6515;
squeal_samples[14590]=8928;
squeal_samples[14591]=11923;
squeal_samples[14592]=14809;
squeal_samples[14593]=17549;
squeal_samples[14594]=20191;
squeal_samples[14595]=22703;
squeal_samples[14596]=25107;
squeal_samples[14597]=27406;
squeal_samples[14598]=29606;
squeal_samples[14599]=31704;
squeal_samples[14600]=33715;
squeal_samples[14601]=35634;
squeal_samples[14602]=37462;
squeal_samples[14603]=39218;
squeal_samples[14604]=40886;
squeal_samples[14605]=42484;
squeal_samples[14606]=44010;
squeal_samples[14607]=45466;
squeal_samples[14608]=46862;
squeal_samples[14609]=48186;
squeal_samples[14610]=49463;
squeal_samples[14611]=50671;
squeal_samples[14612]=51834;
squeal_samples[14613]=52888;
squeal_samples[14614]=49872;
squeal_samples[14615]=44566;
squeal_samples[14616]=39608;
squeal_samples[14617]=34959;
squeal_samples[14618]=30617;
squeal_samples[14619]=26550;
squeal_samples[14620]=22747;
squeal_samples[14621]=19185;
squeal_samples[14622]=15857;
squeal_samples[14623]=12738;
squeal_samples[14624]=9821;
squeal_samples[14625]=7097;
squeal_samples[14626]=7369;
squeal_samples[14627]=10433;
squeal_samples[14628]=13379;
squeal_samples[14629]=16185;
squeal_samples[14630]=18884;
squeal_samples[14631]=21456;
squeal_samples[14632]=23914;
squeal_samples[14633]=26267;
squeal_samples[14634]=28511;
squeal_samples[14635]=30663;
squeal_samples[14636]=32711;
squeal_samples[14637]=34681;
squeal_samples[14638]=36548;
squeal_samples[14639]=38341;
squeal_samples[14640]=40057;
squeal_samples[14641]=41686;
squeal_samples[14642]=43251;
squeal_samples[14643]=44737;
squeal_samples[14644]=46165;
squeal_samples[14645]=47522;
squeal_samples[14646]=48826;
squeal_samples[14647]=50060;
squeal_samples[14648]=51255;
squeal_samples[14649]=52385;
squeal_samples[14650]=52169;
squeal_samples[14651]=47163;
squeal_samples[14652]=42040;
squeal_samples[14653]=37232;
squeal_samples[14654]=32746;
squeal_samples[14655]=28539;
squeal_samples[14656]=24610;
squeal_samples[14657]=20926;
squeal_samples[14658]=17485;
squeal_samples[14659]=14258;
squeal_samples[14660]=11243;
squeal_samples[14661]=8422;
squeal_samples[14662]=6498;
squeal_samples[14663]=8909;
squeal_samples[14664]=11915;
squeal_samples[14665]=14783;
squeal_samples[14666]=17542;
squeal_samples[14667]=20172;
squeal_samples[14668]=22686;
squeal_samples[14669]=25093;
squeal_samples[14670]=27385;
squeal_samples[14671]=29588;
squeal_samples[14672]=31684;
squeal_samples[14673]=33696;
squeal_samples[14674]=35614;
squeal_samples[14675]=37445;
squeal_samples[14676]=39195;
squeal_samples[14677]=40870;
squeal_samples[14678]=42463;
squeal_samples[14679]=43989;
squeal_samples[14680]=45451;
squeal_samples[14681]=46837;
squeal_samples[14682]=48172;
squeal_samples[14683]=49441;
squeal_samples[14684]=50652;
squeal_samples[14685]=51815;
squeal_samples[14686]=52868;
squeal_samples[14687]=49851;
squeal_samples[14688]=44546;
squeal_samples[14689]=39585;
squeal_samples[14690]=34941;
squeal_samples[14691]=30598;
squeal_samples[14692]=26523;
squeal_samples[14693]=22725;
squeal_samples[14694]=19164;
squeal_samples[14695]=15833;
squeal_samples[14696]=12712;
squeal_samples[14697]=9798;
squeal_samples[14698]=7071;
squeal_samples[14699]=7343;
squeal_samples[14700]=10418;
squeal_samples[14701]=13353;
squeal_samples[14702]=16167;
squeal_samples[14703]=18854;
squeal_samples[14704]=21435;
squeal_samples[14705]=23886;
squeal_samples[14706]=26245;
squeal_samples[14707]=28484;
squeal_samples[14708]=30639;
squeal_samples[14709]=32694;
squeal_samples[14710]=34652;
squeal_samples[14711]=36532;
squeal_samples[14712]=38321;
squeal_samples[14713]=40030;
squeal_samples[14714]=41666;
squeal_samples[14715]=43222;
squeal_samples[14716]=44715;
squeal_samples[14717]=46138;
squeal_samples[14718]=47499;
squeal_samples[14719]=48800;
squeal_samples[14720]=50042;
squeal_samples[14721]=51230;
squeal_samples[14722]=52360;
squeal_samples[14723]=52143;
squeal_samples[14724]=47141;
squeal_samples[14725]=42012;
squeal_samples[14726]=37211;
squeal_samples[14727]=32718;
squeal_samples[14728]=28517;
squeal_samples[14729]=24583;
squeal_samples[14730]=20904;
squeal_samples[14731]=17457;
squeal_samples[14732]=14236;
squeal_samples[14733]=11215;
squeal_samples[14734]=8402;
squeal_samples[14735]=6474;
squeal_samples[14736]=8889;
squeal_samples[14737]=11885;
squeal_samples[14738]=14764;
squeal_samples[14739]=17512;
squeal_samples[14740]=20151;
squeal_samples[14741]=22659;
squeal_samples[14742]=25069;
squeal_samples[14743]=27362;
squeal_samples[14744]=29561;
squeal_samples[14745]=31666;
squeal_samples[14746]=33670;
squeal_samples[14747]=35590;
squeal_samples[14748]=37420;
squeal_samples[14749]=39172;
squeal_samples[14750]=40843;
squeal_samples[14751]=42440;
squeal_samples[14752]=43964;
squeal_samples[14753]=45425;
squeal_samples[14754]=46815;
squeal_samples[14755]=48146;
squeal_samples[14756]=49415;
squeal_samples[14757]=50631;
squeal_samples[14758]=51785;
squeal_samples[14759]=52849;
squeal_samples[14760]=49823;
squeal_samples[14761]=44522;
squeal_samples[14762]=39560;
squeal_samples[14763]=34918;
squeal_samples[14764]=30571;
squeal_samples[14765]=26502;
squeal_samples[14766]=22696;
squeal_samples[14767]=19143;
squeal_samples[14768]=15807;
squeal_samples[14769]=12688;
squeal_samples[14770]=9779;
squeal_samples[14771]=7045;
squeal_samples[14772]=7322;
squeal_samples[14773]=10388;
squeal_samples[14774]=13335;
squeal_samples[14775]=16136;
squeal_samples[14776]=18835;
squeal_samples[14777]=21405;
squeal_samples[14778]=23866;
squeal_samples[14779]=26217;
squeal_samples[14780]=28463;
squeal_samples[14781]=30612;
squeal_samples[14782]=32669;
squeal_samples[14783]=34629;
squeal_samples[14784]=36506;
squeal_samples[14785]=38297;
squeal_samples[14786]=40007;
squeal_samples[14787]=41638;
squeal_samples[14788]=43201;
squeal_samples[14789]=44687;
squeal_samples[14790]=46117;
squeal_samples[14791]=47471;
squeal_samples[14792]=48779;
squeal_samples[14793]=50013;
squeal_samples[14794]=51210;
squeal_samples[14795]=52332;
squeal_samples[14796]=52121;
squeal_samples[14797]=47115;
squeal_samples[14798]=41988;
squeal_samples[14799]=37186;
squeal_samples[14800]=32694;
squeal_samples[14801]=28491;
squeal_samples[14802]=24560;
squeal_samples[14803]=20878;
squeal_samples[14804]=17435;
squeal_samples[14805]=14208;
squeal_samples[14806]=11194;
squeal_samples[14807]=8373;
squeal_samples[14808]=6453;
squeal_samples[14809]=8862;
squeal_samples[14810]=11864;
squeal_samples[14811]=14734;
squeal_samples[14812]=17493;
squeal_samples[14813]=20122;
squeal_samples[14814]=22638;
squeal_samples[14815]=25043;
squeal_samples[14816]=27336;
squeal_samples[14817]=29539;
squeal_samples[14818]=31639;
squeal_samples[14819]=33648;
squeal_samples[14820]=35564;
squeal_samples[14821]=37396;
squeal_samples[14822]=39147;
squeal_samples[14823]=40818;
squeal_samples[14824]=42417;
squeal_samples[14825]=43937;
squeal_samples[14826]=45405;
squeal_samples[14827]=46785;
squeal_samples[14828]=48124;
squeal_samples[14829]=49391;
squeal_samples[14830]=50604;
squeal_samples[14831]=51765;
squeal_samples[14832]=52820;
squeal_samples[14833]=49801;
squeal_samples[14834]=44496;
squeal_samples[14835]=39536;
squeal_samples[14836]=34893;
squeal_samples[14837]=30548;
squeal_samples[14838]=26475;
squeal_samples[14839]=22674;
squeal_samples[14840]=19117;
squeal_samples[14841]=15782;
squeal_samples[14842]=12665;
squeal_samples[14843]=9753;
squeal_samples[14844]=7022;
squeal_samples[14845]=7296;
squeal_samples[14846]=10365;
squeal_samples[14847]=13308;
squeal_samples[14848]=16115;
squeal_samples[14849]=18807;
squeal_samples[14850]=21384;
squeal_samples[14851]=23839;
squeal_samples[14852]=26193;
squeal_samples[14853]=28439;
squeal_samples[14854]=30586;
squeal_samples[14855]=32647;
squeal_samples[14856]=34602;
squeal_samples[14857]=36483;
squeal_samples[14858]=38273;
squeal_samples[14859]=39980;
squeal_samples[14860]=41617;
squeal_samples[14861]=43173;
squeal_samples[14862]=44665;
squeal_samples[14863]=46091;
squeal_samples[14864]=47449;
squeal_samples[14865]=48750;
squeal_samples[14866]=49995;
squeal_samples[14867]=51178;
squeal_samples[14868]=52315;
squeal_samples[14869]=52091;
squeal_samples[14870]=47092;
squeal_samples[14871]=41965;
squeal_samples[14872]=37159;
squeal_samples[14873]=32673;
squeal_samples[14874]=28463;
squeal_samples[14875]=24538;
squeal_samples[14876]=20851;
squeal_samples[14877]=17412;
squeal_samples[14878]=14184;
squeal_samples[14879]=11168;
squeal_samples[14880]=8350;
squeal_samples[14881]=6427;
squeal_samples[14882]=8839;
squeal_samples[14883]=11838;
squeal_samples[14884]=14712;
squeal_samples[14885]=17465;
squeal_samples[14886]=20101;
squeal_samples[14887]=22611;
squeal_samples[14888]=25020;
squeal_samples[14889]=27312;
squeal_samples[14890]=29512;
squeal_samples[14891]=31619;
squeal_samples[14892]=33619;
squeal_samples[14893]=35542;
squeal_samples[14894]=37370;
squeal_samples[14895]=39123;
squeal_samples[14896]=40794;
squeal_samples[14897]=42391;
squeal_samples[14898]=43914;
squeal_samples[14899]=45377;
squeal_samples[14900]=46765;
squeal_samples[14901]=48095;
squeal_samples[14902]=49369;
squeal_samples[14903]=50577;
squeal_samples[14904]=51741;
squeal_samples[14905]=52848;
squeal_samples[14906]=50593;
squeal_samples[14907]=45236;
squeal_samples[14908]=40229;
squeal_samples[14909]=35537;
squeal_samples[14910]=31145;
squeal_samples[14911]=27041;
squeal_samples[14912]=23193;
squeal_samples[14913]=19607;
squeal_samples[14914]=16233;
squeal_samples[14915]=13093;
squeal_samples[14916]=10144;
squeal_samples[14917]=7392;
squeal_samples[14918]=6979;
squeal_samples[14919]=10025;
squeal_samples[14920]=12970;
squeal_samples[14921]=15798;
squeal_samples[14922]=18501;
squeal_samples[14923]=21091;
squeal_samples[14924]=23561;
squeal_samples[14925]=25924;
squeal_samples[14926]=28180;
squeal_samples[14927]=30342;
squeal_samples[14928]=32402;
squeal_samples[14929]=34373;
squeal_samples[14930]=36257;
squeal_samples[14931]=38057;
squeal_samples[14932]=39780;
squeal_samples[14933]=41416;
squeal_samples[14934]=42986;
squeal_samples[14935]=44484;
squeal_samples[14936]=45917;
squeal_samples[14937]=47286;
squeal_samples[14938]=48588;
squeal_samples[14939]=49839;
squeal_samples[14940]=51030;
squeal_samples[14941]=52166;
squeal_samples[14942]=52786;
squeal_samples[14943]=48545;
squeal_samples[14944]=43324;
squeal_samples[14945]=38435;
squeal_samples[14946]=33856;
squeal_samples[14947]=29577;
squeal_samples[14948]=25569;
squeal_samples[14949]=21824;
squeal_samples[14950]=18312;
squeal_samples[14951]=15030;
squeal_samples[14952]=11960;
squeal_samples[14953]=9083;
squeal_samples[14954]=6582;
squeal_samples[14955]=8101;
squeal_samples[14956]=11144;
squeal_samples[14957]=14039;
squeal_samples[14958]=16823;
squeal_samples[14959]=19482;
squeal_samples[14960]=22025;
squeal_samples[14961]=24454;
squeal_samples[14962]=26776;
squeal_samples[14963]=28992;
squeal_samples[14964]=31116;
squeal_samples[14965]=33146;
squeal_samples[14966]=35081;
squeal_samples[14967]=36940;
squeal_samples[14968]=38702;
squeal_samples[14969]=40396;
squeal_samples[14970]=42007;
squeal_samples[14971]=43550;
squeal_samples[14972]=45018;
squeal_samples[14973]=46428;
squeal_samples[14974]=47772;
squeal_samples[14975]=49055;
squeal_samples[14976]=50284;
squeal_samples[14977]=51451;
squeal_samples[14978]=52576;
squeal_samples[14979]=51767;
squeal_samples[14980]=46540;
squeal_samples[14981]=41442;
squeal_samples[14982]=36675;
squeal_samples[14983]=32208;
squeal_samples[14984]=28034;
squeal_samples[14985]=24129;
squeal_samples[14986]=20469;
squeal_samples[14987]=17048;
squeal_samples[14988]=13843;
squeal_samples[14989]=10850;
squeal_samples[14990]=8051;
squeal_samples[14991]=6537;
squeal_samples[14992]=9249;
squeal_samples[14993]=12228;
squeal_samples[14994]=15091;
squeal_samples[14995]=17818;
squeal_samples[14996]=20438;
squeal_samples[14997]=22940;
squeal_samples[14998]=25322;
squeal_samples[14999]=27609;
squeal_samples[15000]=29789;
squeal_samples[15001]=31882;
squeal_samples[15002]=33868;
squeal_samples[15003]=35780;
squeal_samples[15004]=37596;
squeal_samples[15005]=39337;
squeal_samples[15006]=40998;
squeal_samples[15007]=42579;
squeal_samples[15008]=44099;
squeal_samples[15009]=45544;
squeal_samples[15010]=46929;
squeal_samples[15011]=48251;
squeal_samples[15012]=49508;
squeal_samples[15013]=50719;
squeal_samples[15014]=51868;
squeal_samples[15015]=52920;
squeal_samples[15016]=49884;
squeal_samples[15017]=44577;
squeal_samples[15018]=39605;
squeal_samples[15019]=34951;
squeal_samples[15020]=30600;
squeal_samples[15021]=26523;
squeal_samples[15022]=22716;
squeal_samples[15023]=19147;
squeal_samples[15024]=15810;
squeal_samples[15025]=12683;
squeal_samples[15026]=9769;
squeal_samples[15027]=7031;
squeal_samples[15028]=7305;
squeal_samples[15029]=10369;
squeal_samples[15030]=13309;
squeal_samples[15031]=16109;
squeal_samples[15032]=18806;
squeal_samples[15033]=21372;
squeal_samples[15034]=23835;
squeal_samples[15035]=26181;
squeal_samples[15036]=28423;
squeal_samples[15037]=30580;
squeal_samples[15038]=32624;
squeal_samples[15039]=34587;
squeal_samples[15040]=36459;
squeal_samples[15041]=38243;
squeal_samples[15042]=39955;
squeal_samples[15043]=41585;
squeal_samples[15044]=43147;
squeal_samples[15045]=44634;
squeal_samples[15046]=46064;
squeal_samples[15047]=47414;
squeal_samples[15048]=48718;
squeal_samples[15049]=49952;
squeal_samples[15050]=51142;
squeal_samples[15051]=52270;
squeal_samples[15052]=52524;
squeal_samples[15053]=47838;
squeal_samples[15054]=42665;
squeal_samples[15055]=37809;
squeal_samples[15056]=33279;
squeal_samples[15057]=29022;
squeal_samples[15058]=25053;
squeal_samples[15059]=21332;
squeal_samples[15060]=17858;
squeal_samples[15061]=14598;
squeal_samples[15062]=11555;
squeal_samples[15063]=8707;
squeal_samples[15064]=6441;
squeal_samples[15065]=8459;
squeal_samples[15066]=11470;
squeal_samples[15067]=14366;
squeal_samples[15068]=17126;
squeal_samples[15069]=19773;
squeal_samples[15070]=22296;
squeal_samples[15071]=24719;
squeal_samples[15072]=27018;
squeal_samples[15073]=29230;
squeal_samples[15074]=31339;
squeal_samples[15075]=33358;
squeal_samples[15076]=35287;
squeal_samples[15077]=37122;
squeal_samples[15078]=38885;
squeal_samples[15079]=40565;
squeal_samples[15080]=42167;
squeal_samples[15081]=43702;
squeal_samples[15082]=45169;
squeal_samples[15083]=46562;
squeal_samples[15084]=47901;
squeal_samples[15085]=49176;
squeal_samples[15086]=50392;
squeal_samples[15087]=51565;
squeal_samples[15088]=52673;
squeal_samples[15089]=51196;
squeal_samples[15090]=45843;
squeal_samples[15091]=40794;
squeal_samples[15092]=36059;
squeal_samples[15093]=31639;
squeal_samples[15094]=27489;
squeal_samples[15095]=23622;
squeal_samples[15096]=19992;
squeal_samples[15097]=16599;
squeal_samples[15098]=13421;
squeal_samples[15099]=10455;
squeal_samples[15100]=7677;
squeal_samples[15101]=6670;
squeal_samples[15102]=9593;
squeal_samples[15103]=12557;
squeal_samples[15104]=15399;
squeal_samples[15105]=18123;
squeal_samples[15106]=20717;
squeal_samples[15107]=23212;
squeal_samples[15108]=25576;
squeal_samples[15109]=27852;
squeal_samples[15110]=30017;
squeal_samples[15111]=32101;
squeal_samples[15112]=34076;
squeal_samples[15113]=35976;
squeal_samples[15114]=37779;
squeal_samples[15115]=39511;
squeal_samples[15116]=41163;
squeal_samples[15117]=42738;
squeal_samples[15118]=44247;
squeal_samples[15119]=45686;
squeal_samples[15120]=47063;
squeal_samples[15121]=48370;
squeal_samples[15122]=49627;
squeal_samples[15123]=50826;
squeal_samples[15124]=51971;
squeal_samples[15125]=52860;
squeal_samples[15126]=49170;
squeal_samples[15127]=43899;
squeal_samples[15128]=38972;
squeal_samples[15129]=34354;
squeal_samples[15130]=30039;
squeal_samples[15131]=25996;
squeal_samples[15132]=22220;
squeal_samples[15133]=18682;
squeal_samples[15134]=15370;
squeal_samples[15135]=12274;
squeal_samples[15136]=9378;
squeal_samples[15137]=6713;
squeal_samples[15138]=7659;
squeal_samples[15139]=10710;
squeal_samples[15140]=13628;
squeal_samples[15141]=16419;
squeal_samples[15142]=19097;
squeal_samples[15143]=21653;
squeal_samples[15144]=24097;
squeal_samples[15145]=26431;
squeal_samples[15146]=28662;
squeal_samples[15147]=30799;
squeal_samples[15148]=32841;
squeal_samples[15149]=34789;
squeal_samples[15150]=36650;
squeal_samples[15151]=38430;
squeal_samples[15152]=40130;
squeal_samples[15153]=41749;
squeal_samples[15154]=43301;
squeal_samples[15155]=44778;
squeal_samples[15156]=46199;
squeal_samples[15157]=47549;
squeal_samples[15158]=48836;
squeal_samples[15159]=50072;
squeal_samples[15160]=51249;
squeal_samples[15161]=52379;
squeal_samples[15162]=52146;
squeal_samples[15163]=47144;
squeal_samples[15164]=41998;
squeal_samples[15165]=37199;
squeal_samples[15166]=32688;
squeal_samples[15167]=28480;
squeal_samples[15168]=24540;
squeal_samples[15169]=20854;
squeal_samples[15170]=17400;
squeal_samples[15171]=14175;
squeal_samples[15172]=11151;
squeal_samples[15173]=8331;
squeal_samples[15174]=6393;
squeal_samples[15175]=8808;
squeal_samples[15176]=11805;
squeal_samples[15177]=14681;
squeal_samples[15178]=17427;
squeal_samples[15179]=20059;
squeal_samples[15180]=22566;
squeal_samples[15181]=24973;
squeal_samples[15182]=27264;
squeal_samples[15183]=29463;
squeal_samples[15184]=31566;
squeal_samples[15185]=33563;
squeal_samples[15186]=35486;
squeal_samples[15187]=37314;
squeal_samples[15188]=39066;
squeal_samples[15189]=40733;
squeal_samples[15190]=42328;
squeal_samples[15191]=43849;
squeal_samples[15192]=45307;
squeal_samples[15193]=46695;
squeal_samples[15194]=48026;
squeal_samples[15195]=49297;
squeal_samples[15196]=50511;
squeal_samples[15197]=51667;
squeal_samples[15198]=52776;
squeal_samples[15199]=50515;
squeal_samples[15200]=45163;
squeal_samples[15201]=40147;
squeal_samples[15202]=35457;
squeal_samples[15203]=31065;
squeal_samples[15204]=26957;
squeal_samples[15205]=23117;
squeal_samples[15206]=19523;
squeal_samples[15207]=16153;
squeal_samples[15208]=13007;
squeal_samples[15209]=10058;
squeal_samples[15210]=7306;
squeal_samples[15211]=6894;
squeal_samples[15212]=9936;
squeal_samples[15213]=12886;
squeal_samples[15214]=15711;
squeal_samples[15215]=18415;
squeal_samples[15216]=21001;
squeal_samples[15217]=23474;
squeal_samples[15218]=25832;
squeal_samples[15219]=28090;
squeal_samples[15220]=30247;
squeal_samples[15221]=32314;
squeal_samples[15222]=34285;
squeal_samples[15223]=36172;
squeal_samples[15224]=37965;
squeal_samples[15225]=39687;
squeal_samples[15226]=41327;
squeal_samples[15227]=42892;
squeal_samples[15228]=44394;
squeal_samples[15229]=45824;
squeal_samples[15230]=47195;
squeal_samples[15231]=48496;
squeal_samples[15232]=49743;
squeal_samples[15233]=50937;
squeal_samples[15234]=52074;
squeal_samples[15235]=52956;
squeal_samples[15236]=49257;
squeal_samples[15237]=43981;
squeal_samples[15238]=39047;
squeal_samples[15239]=34419;
squeal_samples[15240]=30101;
squeal_samples[15241]=26048;
squeal_samples[15242]=22266;
squeal_samples[15243]=18725;
squeal_samples[15244]=15408;
squeal_samples[15245]=12310;
squeal_samples[15246]=9405;
squeal_samples[15247]=6738;
squeal_samples[15248]=7675;
squeal_samples[15249]=10729;
squeal_samples[15250]=13646;
squeal_samples[15251]=16436;
squeal_samples[15252]=19111;
squeal_samples[15253]=21659;
squeal_samples[15254]=24105;
squeal_samples[15255]=26436;
squeal_samples[15256]=28672;
squeal_samples[15257]=30798;
squeal_samples[15258]=32840;
squeal_samples[15259]=34783;
squeal_samples[15260]=36647;
squeal_samples[15261]=38428;
squeal_samples[15262]=40117;
squeal_samples[15263]=41745;
squeal_samples[15264]=43293;
squeal_samples[15265]=44772;
squeal_samples[15266]=46189;
squeal_samples[15267]=47533;
squeal_samples[15268]=48829;
squeal_samples[15269]=50054;
squeal_samples[15270]=51239;
squeal_samples[15271]=52360;
squeal_samples[15272]=52137;
squeal_samples[15273]=47118;
squeal_samples[15274]=41983;
squeal_samples[15275]=37174;
squeal_samples[15276]=32673;
squeal_samples[15277]=28457;
squeal_samples[15278]=24522;
squeal_samples[15279]=20828;
squeal_samples[15280]=17374;
squeal_samples[15281]=14149;
squeal_samples[15282]=11128;
squeal_samples[15283]=8302;
squeal_samples[15284]=6372;
squeal_samples[15285]=8773;
squeal_samples[15286]=11776;
squeal_samples[15287]=14650;
squeal_samples[15288]=17396;
squeal_samples[15289]=20028;
squeal_samples[15290]=22536;
squeal_samples[15291]=24941;
squeal_samples[15292]=27233;
squeal_samples[15293]=29434;
squeal_samples[15294]=31533;
squeal_samples[15295]=33535;
squeal_samples[15296]=35452;
squeal_samples[15297]=37279;
squeal_samples[15298]=39035;
squeal_samples[15299]=40697;
squeal_samples[15300]=42297;
squeal_samples[15301]=43817;
squeal_samples[15302]=45277;
squeal_samples[15303]=46664;
squeal_samples[15304]=47995;
squeal_samples[15305]=49261;
squeal_samples[15306]=50472;
squeal_samples[15307]=51632;
squeal_samples[15308]=52745;
squeal_samples[15309]=51249;
squeal_samples[15310]=45900;
squeal_samples[15311]=40831;
squeal_samples[15312]=36100;
squeal_samples[15313]=31665;
squeal_samples[15314]=27512;
squeal_samples[15315]=23635;
squeal_samples[15316]=20001;
squeal_samples[15317]=16602;
squeal_samples[15318]=13425;
squeal_samples[15319]=10447;
squeal_samples[15320]=7666;
squeal_samples[15321]=6656;
squeal_samples[15322]=9573;
squeal_samples[15323]=12542;
squeal_samples[15324]=15378;
squeal_samples[15325]=18100;
squeal_samples[15326]=20689;
squeal_samples[15327]=23180;
squeal_samples[15328]=25551;
squeal_samples[15329]=27819;
squeal_samples[15330]=29990;
squeal_samples[15331]=32065;
squeal_samples[15332]=34042;
squeal_samples[15333]=35936;
squeal_samples[15334]=37744;
squeal_samples[15335]=39472;
squeal_samples[15336]=41121;
squeal_samples[15337]=42695;
squeal_samples[15338]=44204;
squeal_samples[15339]=45637;
squeal_samples[15340]=47013;
squeal_samples[15341]=48321;
squeal_samples[15342]=49584;
squeal_samples[15343]=50774;
squeal_samples[15344]=51919;
squeal_samples[15345]=52963;
squeal_samples[15346]=49920;
squeal_samples[15347]=44606;
squeal_samples[15348]=39619;
squeal_samples[15349]=34963;
squeal_samples[15350]=30599;
squeal_samples[15351]=26518;
squeal_samples[15352]=22703;
squeal_samples[15353]=19134;
squeal_samples[15354]=15784;
squeal_samples[15355]=12659;
squeal_samples[15356]=9728;
squeal_samples[15357]=6995;
squeal_samples[15358]=7259;
squeal_samples[15359]=10324;
squeal_samples[15360]=13253;
squeal_samples[15361]=16068;
squeal_samples[15362]=18749;
squeal_samples[15363]=21323;
squeal_samples[15364]=23773;
squeal_samples[15365]=26120;
squeal_samples[15366]=28365;
squeal_samples[15367]=30513;
squeal_samples[15368]=32553;
squeal_samples[15369]=34519;
squeal_samples[15370]=36384;
squeal_samples[15371]=38177;
squeal_samples[15372]=39879;
squeal_samples[15373]=41513;
squeal_samples[15374]=43068;
squeal_samples[15375]=44560;
squeal_samples[15376]=45980;
squeal_samples[15377]=47333;
squeal_samples[15378]=48635;
squeal_samples[15379]=49871;
squeal_samples[15380]=51060;
squeal_samples[15381]=52187;
squeal_samples[15382]=52800;
squeal_samples[15383]=48550;
squeal_samples[15384]=43321;
squeal_samples[15385]=38420;
squeal_samples[15386]=33835;
squeal_samples[15387]=29546;
squeal_samples[15388]=25527;
squeal_samples[15389]=21775;
squeal_samples[15390]=18262;
squeal_samples[15391]=14970;
squeal_samples[15392]=11895;
squeal_samples[15393]=9022;
squeal_samples[15394]=6503;
squeal_samples[15395]=8026;
squeal_samples[15396]=11060;
squeal_samples[15397]=13960;
squeal_samples[15398]=16738;
squeal_samples[15399]=19391;
squeal_samples[15400]=21934;
squeal_samples[15401]=24363;
squeal_samples[15402]=26679;
squeal_samples[15403]=28896;
squeal_samples[15404]=31020;
squeal_samples[15405]=33043;
squeal_samples[15406]=34981;
squeal_samples[15407]=36831;
squeal_samples[15408]=38596;
squeal_samples[15409]=40283;
squeal_samples[15410]=41894;
squeal_samples[15411]=43438;
squeal_samples[15412]=44904;
squeal_samples[15413]=46316;
squeal_samples[15414]=47653;
squeal_samples[15415]=48939;
squeal_samples[15416]=50162;
squeal_samples[15417]=51337;
squeal_samples[15418]=52446;
squeal_samples[15419]=52220;
squeal_samples[15420]=47195;
squeal_samples[15421]=42053;
squeal_samples[15422]=37235;
squeal_samples[15423]=32720;
squeal_samples[15424]=28503;
squeal_samples[15425]=24560;
squeal_samples[15426]=20865;
squeal_samples[15427]=17409;
squeal_samples[15428]=14170;
squeal_samples[15429]=11144;
squeal_samples[15430]=8321;
squeal_samples[15431]=6379;
squeal_samples[15432]=8789;
squeal_samples[15433]=11780;
squeal_samples[15434]=14655;
squeal_samples[15435]=17398;
squeal_samples[15436]=20026;
squeal_samples[15437]=22539;
squeal_samples[15438]=24935;
squeal_samples[15439]=27228;
squeal_samples[15440]=29429;
squeal_samples[15441]=31522;
squeal_samples[15442]=33526;
squeal_samples[15443]=35441;
squeal_samples[15444]=37268;
squeal_samples[15445]=39019;
squeal_samples[15446]=40682;
squeal_samples[15447]=42281;
squeal_samples[15448]=43797;
squeal_samples[15449]=45254;
squeal_samples[15450]=46642;
squeal_samples[15451]=47970;
squeal_samples[15452]=49239;
squeal_samples[15453]=50447;
squeal_samples[15454]=51604;
squeal_samples[15455]=52711;
squeal_samples[15456]=51225;
squeal_samples[15457]=45866;
squeal_samples[15458]=40801;
squeal_samples[15459]=36066;
squeal_samples[15460]=31628;
squeal_samples[15461]=27480;
squeal_samples[15462]=23603;
squeal_samples[15463]=19963;
squeal_samples[15464]=16566;
squeal_samples[15465]=13386;
squeal_samples[15466]=10411;
squeal_samples[15467]=7626;
squeal_samples[15468]=6621;
squeal_samples[15469]=9535;
squeal_samples[15470]=12503;
squeal_samples[15471]=15338;
squeal_samples[15472]=18053;
squeal_samples[15473]=20656;
squeal_samples[15474]=23135;
squeal_samples[15475]=25507;
squeal_samples[15476]=27777;
squeal_samples[15477]=29948;
squeal_samples[15478]=32019;
squeal_samples[15479]=34005;
squeal_samples[15480]=35887;
squeal_samples[15481]=37704;
squeal_samples[15482]=39428;
squeal_samples[15483]=41079;
squeal_samples[15484]=42651;
squeal_samples[15485]=44157;
squeal_samples[15486]=45593;
squeal_samples[15487]=46968;
squeal_samples[15488]=48283;
squeal_samples[15489]=49531;
squeal_samples[15490]=50728;
squeal_samples[15491]=51876;
squeal_samples[15492]=52917;
squeal_samples[15493]=49877;
squeal_samples[15494]=44552;
squeal_samples[15495]=39581;
squeal_samples[15496]=34916;
squeal_samples[15497]=30559;
squeal_samples[15498]=26473;
squeal_samples[15499]=22657;
squeal_samples[15500]=19083;
squeal_samples[15501]=15738;
squeal_samples[15502]=12609;
squeal_samples[15503]=9685;
squeal_samples[15504]=6947;
squeal_samples[15505]=7211;
squeal_samples[15506]=10281;
squeal_samples[15507]=13205;
squeal_samples[15508]=16018;
squeal_samples[15509]=18702;
squeal_samples[15510]=21274;
squeal_samples[15511]=23731;
squeal_samples[15512]=26070;
squeal_samples[15513]=28320;
squeal_samples[15514]=30460;
squeal_samples[15515]=32515;
squeal_samples[15516]=34466;
squeal_samples[15517]=36340;
squeal_samples[15518]=38124;
squeal_samples[15519]=39836;
squeal_samples[15520]=41465;
squeal_samples[15521]=43028;
squeal_samples[15522]=44511;
squeal_samples[15523]=45930;
squeal_samples[15524]=47288;
squeal_samples[15525]=48584;
squeal_samples[15526]=49825;
squeal_samples[15527]=51008;
squeal_samples[15528]=52142;
squeal_samples[15529]=52750;
squeal_samples[15530]=48504;
squeal_samples[15531]=43270;
squeal_samples[15532]=38372;
squeal_samples[15533]=33787;
squeal_samples[15534]=29497;
squeal_samples[15535]=25481;
squeal_samples[15536]=21723;
squeal_samples[15537]=18217;
squeal_samples[15538]=14918;
squeal_samples[15539]=11849;
squeal_samples[15540]=8974;
squeal_samples[15541]=6452;
squeal_samples[15542]=7981;
squeal_samples[15543]=11008;
squeal_samples[15544]=13914;
squeal_samples[15545]=16689;
squeal_samples[15546]=19342;
squeal_samples[15547]=21886;
squeal_samples[15548]=24314;
squeal_samples[15549]=26631;
squeal_samples[15550]=28847;
squeal_samples[15551]=30973;
squeal_samples[15552]=32992;
squeal_samples[15553]=34936;
squeal_samples[15554]=36780;
squeal_samples[15555]=38548;
squeal_samples[15556]=40234;
squeal_samples[15557]=41846;
squeal_samples[15558]=43389;
squeal_samples[15559]=44857;
squeal_samples[15560]=46266;
squeal_samples[15561]=47605;
squeal_samples[15562]=48888;
squeal_samples[15563]=50116;
squeal_samples[15564]=51285;
squeal_samples[15565]=52401;
squeal_samples[15566]=52635;
squeal_samples[15567]=47935;
squeal_samples[15568]=42744;
squeal_samples[15569]=37875;
squeal_samples[15570]=33324;
squeal_samples[15571]=29063;
squeal_samples[15572]=25073;
squeal_samples[15573]=21348;
squeal_samples[15574]=17850;
squeal_samples[15575]=14591;
squeal_samples[15576]=11531;
squeal_samples[15577]=8671;
squeal_samples[15578]=6406;
squeal_samples[15579]=8410;
squeal_samples[15580]=11423;
squeal_samples[15581]=14304;
squeal_samples[15582]=17059;
squeal_samples[15583]=19703;
squeal_samples[15584]=22222;
squeal_samples[15585]=24645;
squeal_samples[15586]=26938;
squeal_samples[15587]=29149;
squeal_samples[15588]=31249;
squeal_samples[15589]=33268;
squeal_samples[15590]=35189;
squeal_samples[15591]=37028;
squeal_samples[15592]=38782;
squeal_samples[15593]=40463;
squeal_samples[15594]=42061;
squeal_samples[15595]=43593;
squeal_samples[15596]=45054;
squeal_samples[15597]=46446;
squeal_samples[15598]=47787;
squeal_samples[15599]=49051;
squeal_samples[15600]=50277;
squeal_samples[15601]=51433;
squeal_samples[15602]=52552;
squeal_samples[15603]=51731;
squeal_samples[15604]=46495;
squeal_samples[15605]=41384;
squeal_samples[15606]=36614;
squeal_samples[15607]=32130;
squeal_samples[15608]=27949;
squeal_samples[15609]=24037;
squeal_samples[15610]=20370;
squeal_samples[15611]=16942;
squeal_samples[15612]=13733;
squeal_samples[15613]=10733;
squeal_samples[15614]=7924;
squeal_samples[15615]=6411;
squeal_samples[15616]=9114;
squeal_samples[15617]=12099;
squeal_samples[15618]=14944;
squeal_samples[15619]=17683;
squeal_samples[15620]=20287;
squeal_samples[15621]=22791;
squeal_samples[15622]=25171;
squeal_samples[15623]=27454;
squeal_samples[15624]=29644;
squeal_samples[15625]=31716;
squeal_samples[15626]=33720;
squeal_samples[15627]=35614;
squeal_samples[15628]=37440;
squeal_samples[15629]=39172;
squeal_samples[15630]=40830;
squeal_samples[15631]=42413;
squeal_samples[15632]=43928;
squeal_samples[15633]=45371;
squeal_samples[15634]=46757;
squeal_samples[15635]=48075;
squeal_samples[15636]=49337;
squeal_samples[15637]=50537;
squeal_samples[15638]=51690;
squeal_samples[15639]=52793;
squeal_samples[15640]=51292;
squeal_samples[15641]=45931;
squeal_samples[15642]=40854;
squeal_samples[15643]=36113;
squeal_samples[15644]=31672;
squeal_samples[15645]=27509;
squeal_samples[15646]=23631;
squeal_samples[15647]=19982;
squeal_samples[15648]=16582;
squeal_samples[15649]=13395;
squeal_samples[15650]=10415;
squeal_samples[15651]=7626;
squeal_samples[15652]=6618;
squeal_samples[15653]=9530;
squeal_samples[15654]=12494;
squeal_samples[15655]=15334;
squeal_samples[15656]=18040;
squeal_samples[15657]=20638;
squeal_samples[15658]=23123;
squeal_samples[15659]=25490;
squeal_samples[15660]=27760;
squeal_samples[15661]=29924;
squeal_samples[15662]=31997;
squeal_samples[15663]=33976;
squeal_samples[15664]=35864;
squeal_samples[15665]=37678;
squeal_samples[15666]=39396;
squeal_samples[15667]=41047;
squeal_samples[15668]=42617;
squeal_samples[15669]=44123;
squeal_samples[15670]=45559;
squeal_samples[15671]=46936;
squeal_samples[15672]=48240;
squeal_samples[15673]=49495;
squeal_samples[15674]=50686;
squeal_samples[15675]=51837;
squeal_samples[15676]=52927;
squeal_samples[15677]=50650;
squeal_samples[15678]=45277;
squeal_samples[15679]=40250;
squeal_samples[15680]=35541;
squeal_samples[15681]=31138;
squeal_samples[15682]=27009;
squeal_samples[15683]=23161;
squeal_samples[15684]=19548;
squeal_samples[15685]=16172;
squeal_samples[15686]=13009;
squeal_samples[15687]=10055;
squeal_samples[15688]=7286;
squeal_samples[15689]=6874;
squeal_samples[15690]=9903;
squeal_samples[15691]=12847;
squeal_samples[15692]=15673;
squeal_samples[15693]=18365;
squeal_samples[15694]=20951;
squeal_samples[15695]=23416;
squeal_samples[15696]=25769;
squeal_samples[15697]=28032;
squeal_samples[15698]=30181;
squeal_samples[15699]=32243;
squeal_samples[15700]=34208;
squeal_samples[15701]=36091;
squeal_samples[15702]=37882;
squeal_samples[15703]=39602;
squeal_samples[15704]=41237;
squeal_samples[15705]=42801;
squeal_samples[15706]=44302;
squeal_samples[15707]=45724;
squeal_samples[15708]=47092;
squeal_samples[15709]=48393;
squeal_samples[15710]=49637;
squeal_samples[15711]=50830;
squeal_samples[15712]=51964;
squeal_samples[15713]=52996;
squeal_samples[15714]=49951;
squeal_samples[15715]=44619;
squeal_samples[15716]=39633;
squeal_samples[15717]=34963;
squeal_samples[15718]=30593;
squeal_samples[15719]=26504;
squeal_samples[15720]=22680;
squeal_samples[15721]=19103;
squeal_samples[15722]=15751;
squeal_samples[15723]=12618;
squeal_samples[15724]=9682;
squeal_samples[15725]=6944;
squeal_samples[15726]=7208;
squeal_samples[15727]=10268;
squeal_samples[15728]=13197;
squeal_samples[15729]=16003;
squeal_samples[15730]=18686;
squeal_samples[15731]=21251;
squeal_samples[15732]=23710;
squeal_samples[15733]=26045;
squeal_samples[15734]=28287;
squeal_samples[15735]=30434;
squeal_samples[15736]=32477;
squeal_samples[15737]=34437;
squeal_samples[15738]=36306;
squeal_samples[15739]=38086;
squeal_samples[15740]=39801;
squeal_samples[15741]=41427;
squeal_samples[15742]=42978;
squeal_samples[15743]=44469;
squeal_samples[15744]=45885;
squeal_samples[15745]=47249;
squeal_samples[15746]=48537;
squeal_samples[15747]=49779;
squeal_samples[15748]=50957;
squeal_samples[15749]=52089;
squeal_samples[15750]=52964;
squeal_samples[15751]=49250;
squeal_samples[15752]=43969;
squeal_samples[15753]=39022;
squeal_samples[15754]=34385;
squeal_samples[15755]=30056;
squeal_samples[15756]=25996;
squeal_samples[15757]=22213;
squeal_samples[15758]=18660;
squeal_samples[15759]=15338;
squeal_samples[15760]=12230;
squeal_samples[15761]=9322;
squeal_samples[15762]=6650;
squeal_samples[15763]=7581;
squeal_samples[15764]=10630;
squeal_samples[15765]=13539;
squeal_samples[15766]=16333;
squeal_samples[15767]=18998;
squeal_samples[15768]=21556;
squeal_samples[15769]=23994;
squeal_samples[15770]=26320;
squeal_samples[15771]=28556;
squeal_samples[15772]=30677;
squeal_samples[15773]=32718;
squeal_samples[15774]=34662;
squeal_samples[15775]=36520;
squeal_samples[15776]=38295;
squeal_samples[15777]=39992;
squeal_samples[15778]=41610;
squeal_samples[15779]=43157;
squeal_samples[15780]=44639;
squeal_samples[15781]=46050;
squeal_samples[15782]=47397;
squeal_samples[15783]=48683;
squeal_samples[15784]=49919;
squeal_samples[15785]=51091;
squeal_samples[15786]=52214;
squeal_samples[15787]=52820;
squeal_samples[15788]=48559;
squeal_samples[15789]=43318;
squeal_samples[15790]=38408;
squeal_samples[15791]=33823;
squeal_samples[15792]=29519;
squeal_samples[15793]=25501;
squeal_samples[15794]=21741;
squeal_samples[15795]=18217;
squeal_samples[15796]=14924;
squeal_samples[15797]=11843;
squeal_samples[15798]=8958;
squeal_samples[15799]=6439;
squeal_samples[15800]=7964;
squeal_samples[15801]=10983;
squeal_samples[15802]=13888;
squeal_samples[15803]=16662;
squeal_samples[15804]=19312;
squeal_samples[15805]=21853;
squeal_samples[15806]=24280;
squeal_samples[15807]=26591;
squeal_samples[15808]=28813;
squeal_samples[15809]=30928;
squeal_samples[15810]=32952;
squeal_samples[15811]=34886;
squeal_samples[15812]=36734;
squeal_samples[15813]=38500;
squeal_samples[15814]=40187;
squeal_samples[15815]=41797;
squeal_samples[15816]=43336;
squeal_samples[15817]=44805;
squeal_samples[15818]=46206;
squeal_samples[15819]=47547;
squeal_samples[15820]=48830;
squeal_samples[15821]=50052;
squeal_samples[15822]=51220;
squeal_samples[15823]=52345;
squeal_samples[15824]=52567;
squeal_samples[15825]=47874;
squeal_samples[15826]=42675;
squeal_samples[15827]=37808;
squeal_samples[15828]=33259;
squeal_samples[15829]=28988;
squeal_samples[15830]=25004;
squeal_samples[15831]=21273;
squeal_samples[15832]=17785;
squeal_samples[15833]=14514;
squeal_samples[15834]=11455;
squeal_samples[15835]=8599;
squeal_samples[15836]=6327;
squeal_samples[15837]=8334;
squeal_samples[15838]=11340;
squeal_samples[15839]=14229;
squeal_samples[15840]=16985;
squeal_samples[15841]=19627;
squeal_samples[15842]=22149;
squeal_samples[15843]=24561;
squeal_samples[15844]=26861;
squeal_samples[15845]=29067;
squeal_samples[15846]=31174;
squeal_samples[15847]=33194;
squeal_samples[15848]=35107;
squeal_samples[15849]=36949;
squeal_samples[15850]=38701;
squeal_samples[15851]=40382;
squeal_samples[15852]=41981;
squeal_samples[15853]=43514;
squeal_samples[15854]=44970;
squeal_samples[15855]=46369;
squeal_samples[15856]=47697;
squeal_samples[15857]=48975;
squeal_samples[15858]=50192;
squeal_samples[15859]=51350;
squeal_samples[15860]=52467;
squeal_samples[15861]=52220;
squeal_samples[15862]=47193;
squeal_samples[15863]=42035;
squeal_samples[15864]=37213;
squeal_samples[15865]=32695;
squeal_samples[15866]=28462;
squeal_samples[15867]=24519;
squeal_samples[15868]=20809;
squeal_samples[15869]=17351;
squeal_samples[15870]=14107;
squeal_samples[15871]=11082;
squeal_samples[15872]=8243;
squeal_samples[15873]=6305;
squeal_samples[15874]=8705;
squeal_samples[15875]=11700;
squeal_samples[15876]=14567;
squeal_samples[15877]=17313;
squeal_samples[15878]=19931;
squeal_samples[15879]=22449;
squeal_samples[15880]=24839;
squeal_samples[15881]=27135;
squeal_samples[15882]=29321;
squeal_samples[15883]=31422;
squeal_samples[15884]=33420;
squeal_samples[15885]=35332;
squeal_samples[15886]=37163;
squeal_samples[15887]=38901;
squeal_samples[15888]=40570;
squeal_samples[15889]=42164;
squeal_samples[15890]=43684;
squeal_samples[15891]=45139;
squeal_samples[15892]=46524;
squeal_samples[15893]=47847;
squeal_samples[15894]=49116;
squeal_samples[15895]=50324;
squeal_samples[15896]=51486;
squeal_samples[15897]=52582;
squeal_samples[15898]=52341;
squeal_samples[15899]=47297;
squeal_samples[15900]=42139;
squeal_samples[15901]=37303;
squeal_samples[15902]=32778;
squeal_samples[15903]=28546;
squeal_samples[15904]=24587;
squeal_samples[15905]=20885;
squeal_samples[15906]=17408;
squeal_samples[15907]=14170;
squeal_samples[15908]=11132;
squeal_samples[15909]=8295;
squeal_samples[15910]=6349;
squeal_samples[15911]=8745;
squeal_samples[15912]=11743;
squeal_samples[15913]=14602;
squeal_samples[15914]=17351;
squeal_samples[15915]=19965;
squeal_samples[15916]=22484;
squeal_samples[15917]=24860;
squeal_samples[15918]=27169;
squeal_samples[15919]=29345;
squeal_samples[15920]=31449;
squeal_samples[15921]=33439;
squeal_samples[15922]=35355;
squeal_samples[15923]=37178;
squeal_samples[15924]=38925;
squeal_samples[15925]=40589;
squeal_samples[15926]=42178;
squeal_samples[15927]=43702;
squeal_samples[15928]=45145;
squeal_samples[15929]=46540;
squeal_samples[15930]=47863;
squeal_samples[15931]=49128;
squeal_samples[15932]=50337;
squeal_samples[15933]=51487;
squeal_samples[15934]=52596;
squeal_samples[15935]=51771;
squeal_samples[15936]=46520;
squeal_samples[15937]=41411;
squeal_samples[15938]=36614;
squeal_samples[15939]=32140;
squeal_samples[15940]=27943;
squeal_samples[15941]=24024;
squeal_samples[15942]=20354;
squeal_samples[15943]=16921;
squeal_samples[15944]=13705;
squeal_samples[15945]=10697;
squeal_samples[15946]=7885;
squeal_samples[15947]=6368;
squeal_samples[15948]=9072;
squeal_samples[15949]=12050;
squeal_samples[15950]=14895;
squeal_samples[15951]=17630;
squeal_samples[15952]=20232;
squeal_samples[15953]=22734;
squeal_samples[15954]=25113;
squeal_samples[15955]=27396;
squeal_samples[15956]=29569;
squeal_samples[15957]=31657;
squeal_samples[15958]=33646;
squeal_samples[15959]=35546;
squeal_samples[15960]=37364;
squeal_samples[15961]=39094;
squeal_samples[15962]=40757;
squeal_samples[15963]=42334;
squeal_samples[15964]=43851;
squeal_samples[15965]=45291;
squeal_samples[15966]=46674;
squeal_samples[15967]=47990;
squeal_samples[15968]=49248;
squeal_samples[15969]=50452;
squeal_samples[15970]=51601;
squeal_samples[15971]=52703;
squeal_samples[15972]=51871;
squeal_samples[15973]=46613;
squeal_samples[15974]=41492;
squeal_samples[15975]=36697;
squeal_samples[15976]=32214;
squeal_samples[15977]=28009;
squeal_samples[15978]=24092;
squeal_samples[15979]=20407;
squeal_samples[15980]=16977;
squeal_samples[15981]=13751;
squeal_samples[15982]=10744;
squeal_samples[15983]=7927;
squeal_samples[15984]=6405;
squeal_samples[15985]=9102;
squeal_samples[15986]=12081;
squeal_samples[15987]=14932;
squeal_samples[15988]=17660;
squeal_samples[15989]=20264;
squeal_samples[15990]=22758;
squeal_samples[15991]=25135;
squeal_samples[15992]=27414;
squeal_samples[15993]=29591;
squeal_samples[15994]=31676;
squeal_samples[15995]=33659;
squeal_samples[15996]=35564;
squeal_samples[15997]=37375;
squeal_samples[15998]=39113;
squeal_samples[15999]=40763;
squeal_samples[16000]=42349;
squeal_samples[16001]=43861;
squeal_samples[16002]=45300;
squeal_samples[16003]=46683;
squeal_samples[16004]=47995;
squeal_samples[16005]=49255;
squeal_samples[16006]=50458;
squeal_samples[16007]=51604;
squeal_samples[16008]=52705;
squeal_samples[16009]=51879;
squeal_samples[16010]=46612;
squeal_samples[16011]=41495;
squeal_samples[16012]=36697;
squeal_samples[16013]=32213;
squeal_samples[16014]=28011;
squeal_samples[16015]=24085;
squeal_samples[16016]=20412;
squeal_samples[16017]=16962;
squeal_samples[16018]=13756;
squeal_samples[16019]=10733;
squeal_samples[16020]=7921;
squeal_samples[16021]=6398;
squeal_samples[16022]=9100;
squeal_samples[16023]=12075;
squeal_samples[16024]=14924;
squeal_samples[16025]=17653;
squeal_samples[16026]=20256;
squeal_samples[16027]=22753;
squeal_samples[16028]=25126;
squeal_samples[16029]=27408;
squeal_samples[16030]=29584;
squeal_samples[16031]=31668;
squeal_samples[16032]=33654;
squeal_samples[16033]=35554;
squeal_samples[16034]=37370;
squeal_samples[16035]=39104;
squeal_samples[16036]=40758;
squeal_samples[16037]=42336;
squeal_samples[16038]=43853;
squeal_samples[16039]=45293;
squeal_samples[16040]=46676;
squeal_samples[16041]=47989;
squeal_samples[16042]=49241;
squeal_samples[16043]=50453;
squeal_samples[16044]=51594;
squeal_samples[16045]=52696;
squeal_samples[16046]=51863;
squeal_samples[16047]=46608;
squeal_samples[16048]=41485;
squeal_samples[16049]=36688;
squeal_samples[16050]=32203;
squeal_samples[16051]=27999;
squeal_samples[16052]=24080;
squeal_samples[16053]=20395;
squeal_samples[16054]=16961;
squeal_samples[16055]=13737;
squeal_samples[16056]=10730;
squeal_samples[16057]=7914;
squeal_samples[16058]=6389;
squeal_samples[16059]=9090;
squeal_samples[16060]=12064;
squeal_samples[16061]=14915;
squeal_samples[16062]=17638;
squeal_samples[16063]=20247;
squeal_samples[16064]=22736;
squeal_samples[16065]=25117;
squeal_samples[16066]=27393;
squeal_samples[16067]=29573;
squeal_samples[16068]=31654;
squeal_samples[16069]=33642;
squeal_samples[16070]=35541;
squeal_samples[16071]=37360;
squeal_samples[16072]=39088;
squeal_samples[16073]=40748;
squeal_samples[16074]=42327;
squeal_samples[16075]=43841;
squeal_samples[16076]=45282;
squeal_samples[16077]=46662;
squeal_samples[16078]=47976;
squeal_samples[16079]=49236;
squeal_samples[16080]=50438;
squeal_samples[16081]=51584;
squeal_samples[16082]=52682;
squeal_samples[16083]=51850;
squeal_samples[16084]=46596;
squeal_samples[16085]=41473;
squeal_samples[16086]=36675;
squeal_samples[16087]=32191;
squeal_samples[16088]=27987;
squeal_samples[16089]=24065;
squeal_samples[16090]=20385;
squeal_samples[16091]=16948;
squeal_samples[16092]=13724;
squeal_samples[16093]=10719;
squeal_samples[16094]=7898;
squeal_samples[16095]=6380;
squeal_samples[16096]=9075;
squeal_samples[16097]=12054;
squeal_samples[16098]=14900;
squeal_samples[16099]=17626;
squeal_samples[16100]=20235;
squeal_samples[16101]=22723;
squeal_samples[16102]=25111;
squeal_samples[16103]=27379;
squeal_samples[16104]=29561;
squeal_samples[16105]=31642;
squeal_samples[16106]=33630;
squeal_samples[16107]=35528;
squeal_samples[16108]=37346;
squeal_samples[16109]=39078;
squeal_samples[16110]=40732;
squeal_samples[16111]=42319;
squeal_samples[16112]=43826;
squeal_samples[16113]=45269;
squeal_samples[16114]=46650;
squeal_samples[16115]=47964;
squeal_samples[16116]=49222;
squeal_samples[16117]=50427;
squeal_samples[16118]=51570;
squeal_samples[16119]=52670;
squeal_samples[16120]=51838;
squeal_samples[16121]=46584;
squeal_samples[16122]=41459;
squeal_samples[16123]=36663;
squeal_samples[16124]=32179;
squeal_samples[16125]=27971;
squeal_samples[16126]=24059;
squeal_samples[16127]=20366;
squeal_samples[16128]=16940;
squeal_samples[16129]=13709;
squeal_samples[16130]=10706;
squeal_samples[16131]=7889;
squeal_samples[16132]=6364;
squeal_samples[16133]=9065;
squeal_samples[16134]=12038;
squeal_samples[16135]=14892;
squeal_samples[16136]=17611;
squeal_samples[16137]=20224;
squeal_samples[16138]=22709;
squeal_samples[16139]=25098;
squeal_samples[16140]=27368;
squeal_samples[16141]=29549;
squeal_samples[16142]=31628;
squeal_samples[16143]=33618;
squeal_samples[16144]=35515;
squeal_samples[16145]=37334;
squeal_samples[16146]=39065;
squeal_samples[16147]=40720;
squeal_samples[16148]=42306;
squeal_samples[16149]=43813;
squeal_samples[16150]=45258;
squeal_samples[16151]=46636;
squeal_samples[16152]=47951;
squeal_samples[16153]=49211;
squeal_samples[16154]=50414;
squeal_samples[16155]=51557;
squeal_samples[16156]=52658;
squeal_samples[16157]=51824;
squeal_samples[16158]=46572;
squeal_samples[16159]=41447;
squeal_samples[16160]=36650;
squeal_samples[16161]=32166;
squeal_samples[16162]=27961;
squeal_samples[16163]=24042;
squeal_samples[16164]=20358;
squeal_samples[16165]=16923;
squeal_samples[16166]=13700;
squeal_samples[16167]=10692;
squeal_samples[16168]=7876;
squeal_samples[16169]=6352;
squeal_samples[16170]=9051;
squeal_samples[16171]=12028;
squeal_samples[16172]=14877;
squeal_samples[16173]=17600;
squeal_samples[16174]=20209;
squeal_samples[16175]=22699;
squeal_samples[16176]=25084;
squeal_samples[16177]=27357;
squeal_samples[16178]=29533;
squeal_samples[16179]=31619;
squeal_samples[16180]=33602;
squeal_samples[16181]=35506;
squeal_samples[16182]=37318;
squeal_samples[16183]=39056;
squeal_samples[16184]=40704;
squeal_samples[16185]=42296;
squeal_samples[16186]=43798;
squeal_samples[16187]=45247;
squeal_samples[16188]=46624;
squeal_samples[16189]=47937;
squeal_samples[16190]=49200;
squeal_samples[16191]=50398;
squeal_samples[16192]=51550;
squeal_samples[16193]=52639;
squeal_samples[16194]=51818;
squeal_samples[16195]=46554;
squeal_samples[16196]=41438;
squeal_samples[16197]=36636;
squeal_samples[16198]=32153;
squeal_samples[16199]=27949;
squeal_samples[16200]=24028;
squeal_samples[16201]=20348;
squeal_samples[16202]=16908;
squeal_samples[16203]=13689;
squeal_samples[16204]=10678;
squeal_samples[16205]=7864;
squeal_samples[16206]=6339;
squeal_samples[16207]=9040;
squeal_samples[16208]=12013;
squeal_samples[16209]=14866;
squeal_samples[16210]=17586;
squeal_samples[16211]=20197;
squeal_samples[16212]=22687;
squeal_samples[16213]=25070;
squeal_samples[16214]=27345;
squeal_samples[16215]=29521;
squeal_samples[16216]=31604;
squeal_samples[16217]=33592;
squeal_samples[16218]=35490;
squeal_samples[16219]=37309;
squeal_samples[16220]=39040;
squeal_samples[16221]=40694;
squeal_samples[16222]=42281;
squeal_samples[16223]=43787;
squeal_samples[16224]=45233;
squeal_samples[16225]=46611;
squeal_samples[16226]=47926;
squeal_samples[16227]=49184;
squeal_samples[16228]=50390;
squeal_samples[16229]=51530;
squeal_samples[16230]=52634;
squeal_samples[16231]=52366;
squeal_samples[16232]=47333;
squeal_samples[16233]=42150;
squeal_samples[16234]=37319;
squeal_samples[16235]=32778;
squeal_samples[16236]=28541;
squeal_samples[16237]=24567;
squeal_samples[16238]=20864;
squeal_samples[16239]=17381;
squeal_samples[16240]=14141;
squeal_samples[16241]=11093;
squeal_samples[16242]=8254;
squeal_samples[16243]=6305;
squeal_samples[16244]=8698;
squeal_samples[16245]=11690;
squeal_samples[16246]=14549;
squeal_samples[16247]=17291;
squeal_samples[16248]=19909;
squeal_samples[16249]=22414;
squeal_samples[16250]=24804;
squeal_samples[16251]=27091;
squeal_samples[16252]=29283;
squeal_samples[16253]=31372;
squeal_samples[16254]=33376;
squeal_samples[16255]=35280;
squeal_samples[16256]=37107;
squeal_samples[16257]=38848;
squeal_samples[16258]=40508;
squeal_samples[16259]=42100;
squeal_samples[16260]=43618;
squeal_samples[16261]=45068;
squeal_samples[16262]=46451;
squeal_samples[16263]=47779;
squeal_samples[16264]=49035;
squeal_samples[16265]=50251;
squeal_samples[16266]=51402;
squeal_samples[16267]=52502;
squeal_samples[16268]=52251;
squeal_samples[16269]=47211;
squeal_samples[16270]=42045;
squeal_samples[16271]=37210;
squeal_samples[16272]=32687;
squeal_samples[16273]=28450;
squeal_samples[16274]=24493;
squeal_samples[16275]=20781;
squeal_samples[16276]=17314;
squeal_samples[16277]=14064;
squeal_samples[16278]=11030;
squeal_samples[16279]=8185;
squeal_samples[16280]=6244;
squeal_samples[16281]=8637;
squeal_samples[16282]=11632;
squeal_samples[16283]=14496;
squeal_samples[16284]=17237;
squeal_samples[16285]=19857;
squeal_samples[16286]=22360;
squeal_samples[16287]=24760;
squeal_samples[16288]=27046;
squeal_samples[16289]=29237;
squeal_samples[16290]=31329;
squeal_samples[16291]=33328;
squeal_samples[16292]=35235;
squeal_samples[16293]=37069;
squeal_samples[16294]=38807;
squeal_samples[16295]=40474;
squeal_samples[16296]=42065;
squeal_samples[16297]=43583;
squeal_samples[16298]=45034;
squeal_samples[16299]=46418;
squeal_samples[16300]=47741;
squeal_samples[16301]=49009;
squeal_samples[16302]=50215;
squeal_samples[16303]=51366;
squeal_samples[16304]=52475;
squeal_samples[16305]=52686;
squeal_samples[16306]=47978;
squeal_samples[16307]=42757;
squeal_samples[16308]=37880;
squeal_samples[16309]=33306;
squeal_samples[16310]=29032;
squeal_samples[16311]=25026;
squeal_samples[16312]=21290;
squeal_samples[16313]=17786;
squeal_samples[16314]=14507;
squeal_samples[16315]=11440;
squeal_samples[16316]=8575;
squeal_samples[16317]=6290;
squeal_samples[16318]=8294;
squeal_samples[16319]=11298;
squeal_samples[16320]=14178;
squeal_samples[16321]=16932;
squeal_samples[16322]=19565;
squeal_samples[16323]=22085;
squeal_samples[16324]=24496;
squeal_samples[16325]=26788;
squeal_samples[16326]=28992;
squeal_samples[16327]=31093;
squeal_samples[16328]=33104;
squeal_samples[16329]=35023;
squeal_samples[16330]=36859;
squeal_samples[16331]=38604;
squeal_samples[16332]=40284;
squeal_samples[16333]=41877;
squeal_samples[16334]=43408;
squeal_samples[16335]=44864;
squeal_samples[16336]=46257;
squeal_samples[16337]=47589;
squeal_samples[16338]=48860;
squeal_samples[16339]=50070;
squeal_samples[16340]=51236;
squeal_samples[16341]=52346;
squeal_samples[16342]=52929;
squeal_samples[16343]=48656;
squeal_samples[16344]=43391;
squeal_samples[16345]=38474;
squeal_samples[16346]=33860;
squeal_samples[16347]=29550;
squeal_samples[16348]=25513;
squeal_samples[16349]=21741;
squeal_samples[16350]=18210;
squeal_samples[16351]=14903;
squeal_samples[16352]=11807;
squeal_samples[16353]=8916;
squeal_samples[16354]=6387;
squeal_samples[16355]=7898;
squeal_samples[16356]=10923;
squeal_samples[16357]=13817;
squeal_samples[16358]=16589;
squeal_samples[16359]=19231;
squeal_samples[16360]=21769;
squeal_samples[16361]=24187;
squeal_samples[16362]=26504;
squeal_samples[16363]=28708;
squeal_samples[16364]=30829;
squeal_samples[16365]=32845;
squeal_samples[16366]=34777;
squeal_samples[16367]=36625;
squeal_samples[16368]=38383;
squeal_samples[16369]=40073;
squeal_samples[16370]=41672;
squeal_samples[16371]=43213;
squeal_samples[16372]=44675;
squeal_samples[16373]=46078;
squeal_samples[16374]=47412;
squeal_samples[16375]=48697;
squeal_samples[16376]=49914;
squeal_samples[16377]=51084;
squeal_samples[16378]=52193;
squeal_samples[16379]=53057;
squeal_samples[16380]=49323;
squeal_samples[16381]=44025;
squeal_samples[16382]=39053;
squeal_samples[16383]=34417;
squeal_samples[16384]=30060;
squeal_samples[16385]=25992;
squeal_samples[16386]=22189;
squeal_samples[16387]=18626;
squeal_samples[16388]=15293;
squeal_samples[16389]=12174;
squeal_samples[16390]=9257;
squeal_samples[16391]=6569;
squeal_samples[16392]=7503;
squeal_samples[16393]=10536;
squeal_samples[16394]=13455;
squeal_samples[16395]=16231;
squeal_samples[16396]=18900;
squeal_samples[16397]=21446;
squeal_samples[16398]=23882;
squeal_samples[16399]=26208;
squeal_samples[16400]=28430;
squeal_samples[16401]=30556;
squeal_samples[16402]=32586;
squeal_samples[16403]=34534;
squeal_samples[16404]=36381;
squeal_samples[16405]=38158;
squeal_samples[16406]=39848;
squeal_samples[16407]=41469;
squeal_samples[16408]=43007;
squeal_samples[16409]=44486;
squeal_samples[16410]=45891;
squeal_samples[16411]=47236;
squeal_samples[16412]=48525;
squeal_samples[16413]=49753;
squeal_samples[16414]=50926;
squeal_samples[16415]=52049;
squeal_samples[16416]=53066;
squeal_samples[16417]=50004;
squeal_samples[16418]=44655;
squeal_samples[16419]=39648;
squeal_samples[16420]=34965;
squeal_samples[16421]=30576;
squeal_samples[16422]=26479;
squeal_samples[16423]=22635;
squeal_samples[16424]=19052;
squeal_samples[16425]=15679;
squeal_samples[16426]=12538;
squeal_samples[16427]=9597;
squeal_samples[16428]=6845;
squeal_samples[16429]=7102;
squeal_samples[16430]=10157;
squeal_samples[16431]=13081;
squeal_samples[16432]=15878;
squeal_samples[16433]=18561;
squeal_samples[16434]=21118;
squeal_samples[16435]=23571;
squeal_samples[16436]=25907;
squeal_samples[16437]=28142;
squeal_samples[16438]=30280;
squeal_samples[16439]=32327;
squeal_samples[16440]=34280;
squeal_samples[16441]=36147;
squeal_samples[16442]=37928;
squeal_samples[16443]=39629;
squeal_samples[16444]=41255;
squeal_samples[16445]=42804;
squeal_samples[16446]=44296;
squeal_samples[16447]=45706;
squeal_samples[16448]=47065;
squeal_samples[16449]=48351;
squeal_samples[16450]=49590;
squeal_samples[16451]=50766;
squeal_samples[16452]=51899;
squeal_samples[16453]=52978;
squeal_samples[16454]=50687;
squeal_samples[16455]=45289;
squeal_samples[16456]=40244;
squeal_samples[16457]=35516;
squeal_samples[16458]=31097;
squeal_samples[16459]=26959;
squeal_samples[16460]=23091;
squeal_samples[16461]=19472;
squeal_samples[16462]=16081;
squeal_samples[16463]=12909;
squeal_samples[16464]=9943;
squeal_samples[16465]=7165;
squeal_samples[16466]=6741;
squeal_samples[16467]=9769;
squeal_samples[16468]=12710;
squeal_samples[16469]=15521;
squeal_samples[16470]=18221;
squeal_samples[16471]=20791;
squeal_samples[16472]=23260;
squeal_samples[16473]=25601;
squeal_samples[16474]=27861;
squeal_samples[16475]=30007;
squeal_samples[16476]=32063;
squeal_samples[16477]=34031;
squeal_samples[16478]=35898;
squeal_samples[16479]=37700;
squeal_samples[16480]=39405;
squeal_samples[16481]=41040;
squeal_samples[16482]=42604;
squeal_samples[16483]=44095;
squeal_samples[16484]=45524;
squeal_samples[16485]=46880;
squeal_samples[16486]=48185;
squeal_samples[16487]=49426;
squeal_samples[16488]=50616;
squeal_samples[16489]=51741;
squeal_samples[16490]=52832;
squeal_samples[16491]=51314;
squeal_samples[16492]=45935;
squeal_samples[16493]=40843;
squeal_samples[16494]=36081;
squeal_samples[16495]=31619;
squeal_samples[16496]=27455;
squeal_samples[16497]=23547;
squeal_samples[16498]=19902;
squeal_samples[16499]=16473;
squeal_samples[16500]=13283;
squeal_samples[16501]=10290;
squeal_samples[16502]=7488;
squeal_samples[16503]=6473;
squeal_samples[16504]=9376;
squeal_samples[16505]=12337;
squeal_samples[16506]=15170;
squeal_samples[16507]=17872;
squeal_samples[16508]=20469;
squeal_samples[16509]=22943;
squeal_samples[16510]=25305;
squeal_samples[16511]=27569;
squeal_samples[16512]=29734;
squeal_samples[16513]=31797;
squeal_samples[16514]=33771;
squeal_samples[16515]=35661;
squeal_samples[16516]=37461;
squeal_samples[16517]=39189;
squeal_samples[16518]=40831;
squeal_samples[16519]=42400;
squeal_samples[16520]=43906;
squeal_samples[16521]=45333;
squeal_samples[16522]=46710;
squeal_samples[16523]=48009;
squeal_samples[16524]=49266;
squeal_samples[16525]=50452;
squeal_samples[16526]=51596;
squeal_samples[16527]=52687;
squeal_samples[16528]=51849;
squeal_samples[16529]=46581;
squeal_samples[16530]=41448;
squeal_samples[16531]=36652;
squeal_samples[16532]=32149;
squeal_samples[16533]=27944;
squeal_samples[16534]=24012;
squeal_samples[16535]=20328;
squeal_samples[16536]=16885;
squeal_samples[16537]=13652;
squeal_samples[16538]=10642;
squeal_samples[16539]=7818;
squeal_samples[16540]=6291;
squeal_samples[16541]=8989;
squeal_samples[16542]=11960;
squeal_samples[16543]=14810;
squeal_samples[16544]=17527;
squeal_samples[16545]=20136;
squeal_samples[16546]=22627;
squeal_samples[16547]=25004;
squeal_samples[16548]=27279;
squeal_samples[16549]=29457;
squeal_samples[16550]=31532;
squeal_samples[16551]=33522;
squeal_samples[16552]=35412;
squeal_samples[16553]=37234;
squeal_samples[16554]=38962;
squeal_samples[16555]=40613;
squeal_samples[16556]=42198;
squeal_samples[16557]=43705;
squeal_samples[16558]=45147;
squeal_samples[16559]=46522;
squeal_samples[16560]=47839;
squeal_samples[16561]=49092;
squeal_samples[16562]=50293;
squeal_samples[16563]=51442;
squeal_samples[16564]=52540;
squeal_samples[16565]=52746;
squeal_samples[16566]=48024;
squeal_samples[16567]=42798;
squeal_samples[16568]=37910;
squeal_samples[16569]=33330;
squeal_samples[16570]=29052;
squeal_samples[16571]=25039;
squeal_samples[16572]=21296;
squeal_samples[16573]=17780;
squeal_samples[16574]=14502;
squeal_samples[16575]=11424;
squeal_samples[16576]=8559;
squeal_samples[16577]=6265;
squeal_samples[16578]=8264;
squeal_samples[16579]=11270;
squeal_samples[16580]=14141;
squeal_samples[16581]=16900;
squeal_samples[16582]=19527;
squeal_samples[16583]=22047;
squeal_samples[16584]=24447;
squeal_samples[16585]=26747;
squeal_samples[16586]=28941;
squeal_samples[16587]=31046;
squeal_samples[16588]=33049;
squeal_samples[16589]=34975;
squeal_samples[16590]=36799;
squeal_samples[16591]=38558;
squeal_samples[16592]=40221;
squeal_samples[16593]=41825;
squeal_samples[16594]=43343;
squeal_samples[16595]=44809;
squeal_samples[16596]=46196;
squeal_samples[16597]=47525;
squeal_samples[16598]=48799;
squeal_samples[16599]=50008;
squeal_samples[16600]=51168;
squeal_samples[16601]=52278;
squeal_samples[16602]=52863;
squeal_samples[16603]=48587;
squeal_samples[16604]=43326;
squeal_samples[16605]=38399;
squeal_samples[16606]=33788;
squeal_samples[16607]=29475;
squeal_samples[16608]=25444;
squeal_samples[16609]=21665;
squeal_samples[16610]=18135;
squeal_samples[16611]=14822;
squeal_samples[16612]=11730;
squeal_samples[16613]=8837;
squeal_samples[16614]=6309;
squeal_samples[16615]=7821;
squeal_samples[16616]=10844;
squeal_samples[16617]=13733;
squeal_samples[16618]=16505;
squeal_samples[16619]=19153;
squeal_samples[16620]=21685;
squeal_samples[16621]=24105;
squeal_samples[16622]=26417;
squeal_samples[16623]=28632;
squeal_samples[16624]=30744;
squeal_samples[16625]=32762;
squeal_samples[16626]=34694;
squeal_samples[16627]=36538;
squeal_samples[16628]=38299;
squeal_samples[16629]=39983;
squeal_samples[16630]=41594;
squeal_samples[16631]=43125;
squeal_samples[16632]=44593;
squeal_samples[16633]=45995;
squeal_samples[16634]=47326;
squeal_samples[16635]=48609;
squeal_samples[16636]=49825;
squeal_samples[16637]=50997;
squeal_samples[16638]=52112;
squeal_samples[16639]=53127;
squeal_samples[16640]=50053;
squeal_samples[16641]=44691;
squeal_samples[16642]=39687;
squeal_samples[16643]=34988;
squeal_samples[16644]=30602;
squeal_samples[16645]=26485;
squeal_samples[16646]=22649;
squeal_samples[16647]=19049;
squeal_samples[16648]=15679;
squeal_samples[16649]=12533;
squeal_samples[16650]=9583;
squeal_samples[16651]=6830;
squeal_samples[16652]=7080;
squeal_samples[16653]=10133;
squeal_samples[16654]=13061;
squeal_samples[16655]=15854;
squeal_samples[16656]=18533;
squeal_samples[16657]=21091;
squeal_samples[16658]=23537;
squeal_samples[16659]=25876;
squeal_samples[16660]=28107;
squeal_samples[16661]=30247;
squeal_samples[16662]=32289;
squeal_samples[16663]=34235;
squeal_samples[16664]=36104;
squeal_samples[16665]=37882;
squeal_samples[16666]=39583;
squeal_samples[16667]=41208;
squeal_samples[16668]=42757;
squeal_samples[16669]=44243;
squeal_samples[16670]=45654;
squeal_samples[16671]=47008;
squeal_samples[16672]=48300;
squeal_samples[16673]=49530;
squeal_samples[16674]=50714;
squeal_samples[16675]=51836;
squeal_samples[16676]=52919;
squeal_samples[16677]=51396;
squeal_samples[16678]=46003;
squeal_samples[16679]=40902;
squeal_samples[16680]=36138;
squeal_samples[16681]=31665;
squeal_samples[16682]=27490;
squeal_samples[16683]=23580;
squeal_samples[16684]=19922;
squeal_samples[16685]=16496;
squeal_samples[16686]=13298;
squeal_samples[16687]=10299;
squeal_samples[16688]=7496;
squeal_samples[16689]=6475;
squeal_samples[16690]=9375;
squeal_samples[16691]=12336;
squeal_samples[16692]=15158;
squeal_samples[16693]=17863;
squeal_samples[16694]=20454;
squeal_samples[16695]=22928;
squeal_samples[16696]=25291;
squeal_samples[16697]=27547;
squeal_samples[16698]=29714;
squeal_samples[16699]=31776;
squeal_samples[16700]=33751;
squeal_samples[16701]=35636;
squeal_samples[16702]=37434;
squeal_samples[16703]=39158;
squeal_samples[16704]=40798;
squeal_samples[16705]=42372;
squeal_samples[16706]=43865;
squeal_samples[16707]=45302;
squeal_samples[16708]=46666;
squeal_samples[16709]=47973;
squeal_samples[16710]=49219;
squeal_samples[16711]=50418;
squeal_samples[16712]=51553;
squeal_samples[16713]=52642;
squeal_samples[16714]=52374;
squeal_samples[16715]=47321;
squeal_samples[16716]=42132;
squeal_samples[16717]=37291;
squeal_samples[16718]=32739;
squeal_samples[16719]=28503;
squeal_samples[16720]=24515;
squeal_samples[16721]=20805;
squeal_samples[16722]=17322;
squeal_samples[16723]=14064;
squeal_samples[16724]=11017;
squeal_samples[16725]=8168;
squeal_samples[16726]=6216;
squeal_samples[16727]=8604;
squeal_samples[16728]=11592;
squeal_samples[16729]=14452;
squeal_samples[16730]=17188;
squeal_samples[16731]=19805;
squeal_samples[16732]=22308;
squeal_samples[16733]=24697;
squeal_samples[16734]=26980;
squeal_samples[16735]=29172;
squeal_samples[16736]=31256;
squeal_samples[16737]=33252;
squeal_samples[16738]=35160;
squeal_samples[16739]=36977;
squeal_samples[16740]=38723;
squeal_samples[16741]=40377;
squeal_samples[16742]=41975;
squeal_samples[16743]=43483;
squeal_samples[16744]=44936;
squeal_samples[16745]=46318;
squeal_samples[16746]=47638;
squeal_samples[16747]=48905;
squeal_samples[16748]=50108;
squeal_samples[16749]=51266;
squeal_samples[16750]=52359;
squeal_samples[16751]=52946;
squeal_samples[16752]=48658;
squeal_samples[16753]=43389;
squeal_samples[16754]=38457;
squeal_samples[16755]=33841;
squeal_samples[16756]=29520;
squeal_samples[16757]=25481;
squeal_samples[16758]=21694;
squeal_samples[16759]=18160;
squeal_samples[16760]=14843;
squeal_samples[16761]=11748;
squeal_samples[16762]=8852;
squeal_samples[16763]=6318;
squeal_samples[16764]=7824;
squeal_samples[16765]=10846;
squeal_samples[16766]=13738;
squeal_samples[16767]=16502;
squeal_samples[16768]=19151;
squeal_samples[16769]=21684;
squeal_samples[16770]=24095;
squeal_samples[16771]=26413;
squeal_samples[16772]=28617;
squeal_samples[16773]=30730;
squeal_samples[16774]=32750;
squeal_samples[16775]=34675;
squeal_samples[16776]=36521;
squeal_samples[16777]=38280;
squeal_samples[16778]=39958;
squeal_samples[16779]=41571;
squeal_samples[16780]=43100;
squeal_samples[16781]=44572;
squeal_samples[16782]=45962;
squeal_samples[16783]=47307;
squeal_samples[16784]=48579;
squeal_samples[16785]=49801;
squeal_samples[16786]=50965;
squeal_samples[16787]=52079;
squeal_samples[16788]=53093;
squeal_samples[16789]=50015;
squeal_samples[16790]=44661;
squeal_samples[16791]=39641;
squeal_samples[16792]=34955;
squeal_samples[16793]=30561;
squeal_samples[16794]=26450;
squeal_samples[16795]=22606;
squeal_samples[16796]=19009;
squeal_samples[16797]=15641;
squeal_samples[16798]=12490;
squeal_samples[16799]=9546;
squeal_samples[16800]=6789;
squeal_samples[16801]=7037;
squeal_samples[16802]=10093;
squeal_samples[16803]=13010;
squeal_samples[16804]=15814;
squeal_samples[16805]=18484;
squeal_samples[16806]=21047;
squeal_samples[16807]=23491;
squeal_samples[16808]=25830;
squeal_samples[16809]=28063;
squeal_samples[16810]=30201;
squeal_samples[16811]=32244;
squeal_samples[16812]=34189;
squeal_samples[16813]=36059;
squeal_samples[16814]=37837;
squeal_samples[16815]=39535;
squeal_samples[16816]=41161;
squeal_samples[16817]=42708;
squeal_samples[16818]=44196;
squeal_samples[16819]=45606;
squeal_samples[16820]=46963;
squeal_samples[16821]=48254;
squeal_samples[16822]=49486;
squeal_samples[16823]=50668;
squeal_samples[16824]=51791;
squeal_samples[16825]=52873;
squeal_samples[16826]=51347;
squeal_samples[16827]=45955;
squeal_samples[16828]=40860;
squeal_samples[16829]=36084;
squeal_samples[16830]=31621;
squeal_samples[16831]=27439;
squeal_samples[16832]=23537;
squeal_samples[16833]=19872;
squeal_samples[16834]=16451;
squeal_samples[16835]=13242;
squeal_samples[16836]=10250;
squeal_samples[16837]=7447;
squeal_samples[16838]=6421;
squeal_samples[16839]=9328;
squeal_samples[16840]=12282;
squeal_samples[16841]=15109;
squeal_samples[16842]=17817;
squeal_samples[16843]=20403;
squeal_samples[16844]=22878;
squeal_samples[16845]=25240;
squeal_samples[16846]=27501;
squeal_samples[16847]=29665;
squeal_samples[16848]=31724;
squeal_samples[16849]=33701;
squeal_samples[16850]=35584;
squeal_samples[16851]=37384;
squeal_samples[16852]=39107;
squeal_samples[16853]=40749;
squeal_samples[16854]=42319;
squeal_samples[16855]=43816;
squeal_samples[16856]=45249;
squeal_samples[16857]=46618;
squeal_samples[16858]=47920;
squeal_samples[16859]=49171;
squeal_samples[16860]=50364;
squeal_samples[16861]=51505;
squeal_samples[16862]=52589;
squeal_samples[16863]=52326;
squeal_samples[16864]=47267;
squeal_samples[16865]=42086;
squeal_samples[16866]=37234;
squeal_samples[16867]=32695;
squeal_samples[16868]=28446;
squeal_samples[16869]=24469;
squeal_samples[16870]=20752;
squeal_samples[16871]=17273;
squeal_samples[16872]=14011;
squeal_samples[16873]=10968;
squeal_samples[16874]=8116;
squeal_samples[16875]=6166;
squeal_samples[16876]=8560;
squeal_samples[16877]=11539;
squeal_samples[16878]=14404;
squeal_samples[16879]=17133;
squeal_samples[16880]=19758;
squeal_samples[16881]=22255;
squeal_samples[16882]=24648;
squeal_samples[16883]=26929;
squeal_samples[16884]=29120;
squeal_samples[16885]=31206;
squeal_samples[16886]=33200;
squeal_samples[16887]=35110;
squeal_samples[16888]=36927;
squeal_samples[16889]=38670;
squeal_samples[16890]=40330;
squeal_samples[16891]=41920;
squeal_samples[16892]=43434;
squeal_samples[16893]=44884;
squeal_samples[16894]=46267;
squeal_samples[16895]=47589;
squeal_samples[16896]=48851;
squeal_samples[16897]=50062;
squeal_samples[16898]=51209;
squeal_samples[16899]=52312;
squeal_samples[16900]=53153;
squeal_samples[16901]=49411;
squeal_samples[16902]=44097;
squeal_samples[16903]=39109;
squeal_samples[16904]=34453;
squeal_samples[16905]=30085;
squeal_samples[16906]=26001;
squeal_samples[16907]=22192;
squeal_samples[16908]=18609;
squeal_samples[16909]=15269;
squeal_samples[16910]=12133;
squeal_samples[16911]=9219;
squeal_samples[16912]=6517;
squeal_samples[16913]=7451;
squeal_samples[16914]=10472;
squeal_samples[16915]=13385;
squeal_samples[16916]=16162;
squeal_samples[16917]=18820;
squeal_samples[16918]=21364;
squeal_samples[16919]=23797;
squeal_samples[16920]=26116;
squeal_samples[16921]=28334;
squeal_samples[16922]=30457;
squeal_samples[16923]=32488;
squeal_samples[16924]=34421;
squeal_samples[16925]=36279;
squeal_samples[16926]=38039;
squeal_samples[16927]=39740;
squeal_samples[16928]=41347;
squeal_samples[16929]=42889;
squeal_samples[16930]=44363;
squeal_samples[16931]=45765;
squeal_samples[16932]=47114;
squeal_samples[16933]=48394;
squeal_samples[16934]=49623;
squeal_samples[16935]=50791;
squeal_samples[16936]=51912;
squeal_samples[16937]=52980;
squeal_samples[16938]=51451;
squeal_samples[16939]=46047;
squeal_samples[16940]=40941;
squeal_samples[16941]=36159;
squeal_samples[16942]=31693;
squeal_samples[16943]=27504;
squeal_samples[16944]=23588;
squeal_samples[16945]=19927;
squeal_samples[16946]=16492;
squeal_samples[16947]=13292;
squeal_samples[16948]=10279;
squeal_samples[16949]=7480;
squeal_samples[16950]=6448;
squeal_samples[16951]=9351;
squeal_samples[16952]=12301;
squeal_samples[16953]=15134;
squeal_samples[16954]=17831;
squeal_samples[16955]=20420;
squeal_samples[16956]=22889;
squeal_samples[16957]=25249;
squeal_samples[16958]=27510;
squeal_samples[16959]=29666;
squeal_samples[16960]=31733;
squeal_samples[16961]=33698;
squeal_samples[16962]=35585;
squeal_samples[16963]=37386;
squeal_samples[16964]=39097;
squeal_samples[16965]=40748;
squeal_samples[16966]=42310;
squeal_samples[16967]=43811;
squeal_samples[16968]=45240;
squeal_samples[16969]=46605;
squeal_samples[16970]=47909;
squeal_samples[16971]=49161;
squeal_samples[16972]=50346;
squeal_samples[16973]=51489;
squeal_samples[16974]=52572;
squeal_samples[16975]=52776;
squeal_samples[16976]=48039;
squeal_samples[16977]=42808;
squeal_samples[16978]=37908;
squeal_samples[16979]=33323;
squeal_samples[16980]=29031;
squeal_samples[16981]=25013;
squeal_samples[16982]=21260;
squeal_samples[16983]=17742;
squeal_samples[16984]=14455;
squeal_samples[16985]=11373;
squeal_samples[16986]=8497;
squeal_samples[16987]=6205;
squeal_samples[16988]=8197;
squeal_samples[16989]=11203;
squeal_samples[16990]=14071;
squeal_samples[16991]=16824;
squeal_samples[16992]=19451;
squeal_samples[16993]=21962;
squeal_samples[16994]=24367;
squeal_samples[16995]=26656;
squeal_samples[16996]=28860;
squeal_samples[16997]=30953;
squeal_samples[16998]=32959;
squeal_samples[16999]=34878;
squeal_samples[17000]=36704;
squeal_samples[17001]=38453;
squeal_samples[17002]=40124;
squeal_samples[17003]=41719;
squeal_samples[17004]=43245;
squeal_samples[17005]=44699;
squeal_samples[17006]=46089;
squeal_samples[17007]=47419;
squeal_samples[17008]=48685;
squeal_samples[17009]=49896;
squeal_samples[17010]=51053;
squeal_samples[17011]=52161;
squeal_samples[17012]=53166;
squeal_samples[17013]=50084;
squeal_samples[17014]=44718;
squeal_samples[17015]=39691;
squeal_samples[17016]=34998;
squeal_samples[17017]=30594;
squeal_samples[17018]=26476;
squeal_samples[17019]=22630;
squeal_samples[17020]=19022;
squeal_samples[17021]=15650;
squeal_samples[17022]=12487;
squeal_samples[17023]=9544;
squeal_samples[17024]=6775;
squeal_samples[17025]=7030;
squeal_samples[17026]=10077;
squeal_samples[17027]=13000;
squeal_samples[17028]=15785;
squeal_samples[17029]=18470;
squeal_samples[17030]=21019;
squeal_samples[17031]=23470;
squeal_samples[17032]=25797;
squeal_samples[17033]=28035;
squeal_samples[17034]=30166;
squeal_samples[17035]=32208;
squeal_samples[17036]=34150;
squeal_samples[17037]=36021;
squeal_samples[17038]=37794;
squeal_samples[17039]=39493;
squeal_samples[17040]=41115;
squeal_samples[17041]=42668;
squeal_samples[17042]=44149;
squeal_samples[17043]=45560;
squeal_samples[17044]=46914;
squeal_samples[17045]=48202;
squeal_samples[17046]=49442;
squeal_samples[17047]=50608;
squeal_samples[17048]=51742;
squeal_samples[17049]=52813;
squeal_samples[17050]=51971;
squeal_samples[17051]=46674;
squeal_samples[17052]=41531;
squeal_samples[17053]=36707;
squeal_samples[17054]=32198;
squeal_samples[17055]=27977;
squeal_samples[17056]=24028;
squeal_samples[17057]=20333;
squeal_samples[17058]=16871;
squeal_samples[17059]=13641;
squeal_samples[17060]=10615;
squeal_samples[17061]=7781;
squeal_samples[17062]=6245;
squeal_samples[17063]=8935;
squeal_samples[17064]=11903;
squeal_samples[17065]=14745;
squeal_samples[17066]=17465;
squeal_samples[17067]=20065;
squeal_samples[17068]=22555;
squeal_samples[17069]=24916;
squeal_samples[17070]=27197;
squeal_samples[17071]=29362;
squeal_samples[17072]=31440;
squeal_samples[17073]=33422;
squeal_samples[17074]=35320;
squeal_samples[17075]=37123;
squeal_samples[17076]=38858;
squeal_samples[17077]=40504;
squeal_samples[17078]=42083;
squeal_samples[17079]=43585;
squeal_samples[17080]=45029;
squeal_samples[17081]=46399;
squeal_samples[17082]=47716;
squeal_samples[17083]=48969;
squeal_samples[17084]=50164;
squeal_samples[17085]=51312;
squeal_samples[17086]=52406;
squeal_samples[17087]=52982;
squeal_samples[17088]=48681;
squeal_samples[17089]=43406;
squeal_samples[17090]=38467;
squeal_samples[17091]=33842;
squeal_samples[17092]=29511;
squeal_samples[17093]=25462;
squeal_samples[17094]=21676;
squeal_samples[17095]=18130;
squeal_samples[17096]=14813;
squeal_samples[17097]=11710;
squeal_samples[17098]=8809;
squeal_samples[17099]=6269;
squeal_samples[17100]=7775;
squeal_samples[17101]=10794;
squeal_samples[17102]=13682;
squeal_samples[17103]=16450;
squeal_samples[17104]=19091;
squeal_samples[17105]=21618;
squeal_samples[17106]=24038;
squeal_samples[17107]=26339;
squeal_samples[17108]=28551;
squeal_samples[17109]=30658;
squeal_samples[17110]=32681;
squeal_samples[17111]=34604;
squeal_samples[17112]=36445;
squeal_samples[17113]=38205;
squeal_samples[17114]=39878;
squeal_samples[17115]=41489;
squeal_samples[17116]=43015;
squeal_samples[17117]=44484;
squeal_samples[17118]=45882;
squeal_samples[17119]=47220;
squeal_samples[17120]=48488;
squeal_samples[17121]=49713;
squeal_samples[17122]=50876;
squeal_samples[17123]=51982;
squeal_samples[17124]=53059;
squeal_samples[17125]=50741;
squeal_samples[17126]=45336;
squeal_samples[17127]=40268;
squeal_samples[17128]=35528;
squeal_samples[17129]=31092;
squeal_samples[17130]=26936;
squeal_samples[17131]=23059;
squeal_samples[17132]=19422;
squeal_samples[17133]=16020;
squeal_samples[17134]=12842;
squeal_samples[17135]=9859;
squeal_samples[17136]=7080;
squeal_samples[17137]=6641;
squeal_samples[17138]=9667;
squeal_samples[17139]=12601;
squeal_samples[17140]=15409;
squeal_samples[17141]=18098;
squeal_samples[17142]=20670;
squeal_samples[17143]=23132;
squeal_samples[17144]=25473;
squeal_samples[17145]=27725;
squeal_samples[17146]=29863;
squeal_samples[17147]=31920;
squeal_samples[17148]=33875;
squeal_samples[17149]=35756;
squeal_samples[17150]=37539;
squeal_samples[17151]=39249;
squeal_samples[17152]=40883;
squeal_samples[17153]=42439;
squeal_samples[17154]=43929;
squeal_samples[17155]=45348;
squeal_samples[17156]=46714;
squeal_samples[17157]=48008;
squeal_samples[17158]=49251;
squeal_samples[17159]=50431;
squeal_samples[17160]=51566;
squeal_samples[17161]=52648;
squeal_samples[17162]=52375;
squeal_samples[17163]=47309;
squeal_samples[17164]=42116;
squeal_samples[17165]=37252;
squeal_samples[17166]=32708;
squeal_samples[17167]=28450;
squeal_samples[17168]=24470;
squeal_samples[17169]=20744;
squeal_samples[17170]=17260;
squeal_samples[17171]=13993;
squeal_samples[17172]=10941;
squeal_samples[17173]=8088;
squeal_samples[17174]=6130;
squeal_samples[17175]=8518;
squeal_samples[17176]=11502;
squeal_samples[17177]=14359;
squeal_samples[17178]=17091;
squeal_samples[17179]=19708;
squeal_samples[17180]=22207;
squeal_samples[17181]=24593;
squeal_samples[17182]=26881;
squeal_samples[17183]=29060;
squeal_samples[17184]=31151;
squeal_samples[17185]=33144;
squeal_samples[17186]=35045;
squeal_samples[17187]=36867;
squeal_samples[17188]=38606;
squeal_samples[17189]=40268;
squeal_samples[17190]=41853;
squeal_samples[17191]=43367;
squeal_samples[17192]=44814;
squeal_samples[17193]=46198;
squeal_samples[17194]=47510;
squeal_samples[17195]=48784;
squeal_samples[17196]=49977;
squeal_samples[17197]=51136;
squeal_samples[17198]=52231;
squeal_samples[17199]=53074;
squeal_samples[17200]=49330;
squeal_samples[17201]=44008;
squeal_samples[17202]=39030;
squeal_samples[17203]=34366;
squeal_samples[17204]=30002;
squeal_samples[17205]=25919;
squeal_samples[17206]=22099;
squeal_samples[17207]=18530;
squeal_samples[17208]=15180;
squeal_samples[17209]=12049;
squeal_samples[17210]=9124;
squeal_samples[17211]=6428;
squeal_samples[17212]=7352;
squeal_samples[17213]=10387;
squeal_samples[17214]=13291;
squeal_samples[17215]=16072;
squeal_samples[17216]=18725;
squeal_samples[17217]=21276;
squeal_samples[17218]=23696;
squeal_samples[17219]=26027;
squeal_samples[17220]=28234;
squeal_samples[17221]=30368;
squeal_samples[17222]=32387;
squeal_samples[17223]=34333;
squeal_samples[17224]=36178;
squeal_samples[17225]=37949;
squeal_samples[17226]=39644;
squeal_samples[17227]=41251;
squeal_samples[17228]=42797;
squeal_samples[17229]=44265;
squeal_samples[17230]=45672;
squeal_samples[17231]=47014;
squeal_samples[17232]=48299;
squeal_samples[17233]=49523;
squeal_samples[17234]=50695;
squeal_samples[17235]=51812;
squeal_samples[17236]=52885;
squeal_samples[17237]=52025;
squeal_samples[17238]=46728;
squeal_samples[17239]=41575;
squeal_samples[17240]=36749;
squeal_samples[17241]=32233;
squeal_samples[17242]=28001;
squeal_samples[17243]=24055;
squeal_samples[17244]=20348;
squeal_samples[17245]=16888;
squeal_samples[17246]=13641;
squeal_samples[17247]=10614;
squeal_samples[17248]=7779;
squeal_samples[17249]=6241;
squeal_samples[17250]=8927;
squeal_samples[17251]=11896;
squeal_samples[17252]=14730;
squeal_samples[17253]=17448;
squeal_samples[17254]=20046;
squeal_samples[17255]=22533;
squeal_samples[17256]=24903;
squeal_samples[17257]=27166;
squeal_samples[17258]=29344;
squeal_samples[17259]=31411;
squeal_samples[17260]=33395;
squeal_samples[17261]=35290;
squeal_samples[17262]=37092;
squeal_samples[17263]=38824;
squeal_samples[17264]=40469;
squeal_samples[17265]=42045;
squeal_samples[17266]=43554;
squeal_samples[17267]=44991;
squeal_samples[17268]=46365;
squeal_samples[17269]=47675;
squeal_samples[17270]=48927;
squeal_samples[17271]=50125;
squeal_samples[17272]=51264;
squeal_samples[17273]=52361;
squeal_samples[17274]=53195;
squeal_samples[17275]=49446;
squeal_samples[17276]=44114;
squeal_samples[17277]=39122;
squeal_samples[17278]=34452;
squeal_samples[17279]=30080;
squeal_samples[17280]=25990;
squeal_samples[17281]=22169;
squeal_samples[17282]=18588;
squeal_samples[17283]=15235;
squeal_samples[17284]=12097;
squeal_samples[17285]=9173;
squeal_samples[17286]=6464;
squeal_samples[17287]=7396;
squeal_samples[17288]=10418;
squeal_samples[17289]=13324;
squeal_samples[17290]=16098;
squeal_samples[17291]=18758;
squeal_samples[17292]=21295;
squeal_samples[17293]=23727;
squeal_samples[17294]=26042;
squeal_samples[17295]=28262;
squeal_samples[17296]=30377;
squeal_samples[17297]=32414;
squeal_samples[17298]=34340;
squeal_samples[17299]=36195;
squeal_samples[17300]=37960;
squeal_samples[17301]=39651;
squeal_samples[17302]=41261;
squeal_samples[17303]=42798;
squeal_samples[17304]=44268;
squeal_samples[17305]=45675;
squeal_samples[17306]=47013;
squeal_samples[17307]=48299;
squeal_samples[17308]=49523;
squeal_samples[17309]=50695;
squeal_samples[17310]=51807;
squeal_samples[17311]=52883;
squeal_samples[17312]=52019;
squeal_samples[17313]=46728;
squeal_samples[17314]=41564;
squeal_samples[17315]=36744;
squeal_samples[17316]=32221;
squeal_samples[17317]=27996;
squeal_samples[17318]=24037;
squeal_samples[17319]=20338;
squeal_samples[17320]=16872;
squeal_samples[17321]=13628;
squeal_samples[17322]=10600;
squeal_samples[17323]=7760;
squeal_samples[17324]=6220;
squeal_samples[17325]=8916;
squeal_samples[17326]=11873;
squeal_samples[17327]=14719;
squeal_samples[17328]=17433;
squeal_samples[17329]=20026;
squeal_samples[17330]=22516;
squeal_samples[17331]=24881;
squeal_samples[17332]=27149;
squeal_samples[17333]=29322;
squeal_samples[17334]=31394;
squeal_samples[17335]=33376;
squeal_samples[17336]=35268;
squeal_samples[17337]=37077;
squeal_samples[17338]=38800;
squeal_samples[17339]=40453;
squeal_samples[17340]=42025;
squeal_samples[17341]=43534;
squeal_samples[17342]=44967;
squeal_samples[17343]=46341;
squeal_samples[17344]=47654;
squeal_samples[17345]=48904;
squeal_samples[17346]=50104;
squeal_samples[17347]=51247;
squeal_samples[17348]=52340;
squeal_samples[17349]=53177;
squeal_samples[17350]=49421;
squeal_samples[17351]=44088;
squeal_samples[17352]=39106;
squeal_samples[17353]=34430;
squeal_samples[17354]=30062;
squeal_samples[17355]=25971;
squeal_samples[17356]=22149;
squeal_samples[17357]=18565;
squeal_samples[17358]=15215;
squeal_samples[17359]=12078;
squeal_samples[17360]=9147;
squeal_samples[17361]=6448;
squeal_samples[17362]=7367;
squeal_samples[17363]=10398;
squeal_samples[17364]=13297;
squeal_samples[17365]=16078;
squeal_samples[17366]=18737;
squeal_samples[17367]=21272;
squeal_samples[17368]=23704;
squeal_samples[17369]=26018;
squeal_samples[17370]=28241;
squeal_samples[17371]=30356;
squeal_samples[17372]=32386;
squeal_samples[17373]=34318;
squeal_samples[17374]=36167;
squeal_samples[17375]=37939;
squeal_samples[17376]=39624;
squeal_samples[17377]=41238;
squeal_samples[17378]=42779;
squeal_samples[17379]=44246;
squeal_samples[17380]=45654;
squeal_samples[17381]=46986;
squeal_samples[17382]=48276;
squeal_samples[17383]=49498;
squeal_samples[17384]=50669;
squeal_samples[17385]=51789;
squeal_samples[17386]=52858;
squeal_samples[17387]=51995;
squeal_samples[17388]=46703;
squeal_samples[17389]=41540;
squeal_samples[17390]=36717;
squeal_samples[17391]=32201;
squeal_samples[17392]=27964;
squeal_samples[17393]=24020;
squeal_samples[17394]=20309;
squeal_samples[17395]=16849;
squeal_samples[17396]=13605;
squeal_samples[17397]=10572;
squeal_samples[17398]=7737;
squeal_samples[17399]=6197;
squeal_samples[17400]=8888;
squeal_samples[17401]=11854;
squeal_samples[17402]=14689;
squeal_samples[17403]=17412;
squeal_samples[17404]=19999;
squeal_samples[17405]=22494;
squeal_samples[17406]=24853;
squeal_samples[17407]=27134;
squeal_samples[17408]=29294;
squeal_samples[17409]=31372;
squeal_samples[17410]=33349;
squeal_samples[17411]=35245;
squeal_samples[17412]=37052;
squeal_samples[17413]=38776;
squeal_samples[17414]=40429;
squeal_samples[17415]=41998;
squeal_samples[17416]=43512;
squeal_samples[17417]=44942;
squeal_samples[17418]=46315;
squeal_samples[17419]=47631;
squeal_samples[17420]=48879;
squeal_samples[17421]=50080;
squeal_samples[17422]=51222;
squeal_samples[17423]=52316;
squeal_samples[17424]=53151;
squeal_samples[17425]=49397;
squeal_samples[17426]=44065;
squeal_samples[17427]=39080;
squeal_samples[17428]=34405;
squeal_samples[17429]=30039;
squeal_samples[17430]=25944;
squeal_samples[17431]=22128;
squeal_samples[17432]=18537;
squeal_samples[17433]=15192;
squeal_samples[17434]=12053;
squeal_samples[17435]=9122;
squeal_samples[17436]=6425;
squeal_samples[17437]=7342;
squeal_samples[17438]=10372;
squeal_samples[17439]=13274;
squeal_samples[17440]=16053;
squeal_samples[17441]=18711;
squeal_samples[17442]=21250;
squeal_samples[17443]=23677;
squeal_samples[17444]=25996;
squeal_samples[17445]=28214;
squeal_samples[17446]=30333;
squeal_samples[17447]=32360;
squeal_samples[17448]=34295;
squeal_samples[17449]=36143;
squeal_samples[17450]=37913;
squeal_samples[17451]=39601;
squeal_samples[17452]=41212;
squeal_samples[17453]=42754;
squeal_samples[17454]=44225;
squeal_samples[17455]=45625;
squeal_samples[17456]=46966;
squeal_samples[17457]=48248;
squeal_samples[17458]=49474;
squeal_samples[17459]=50647;
squeal_samples[17460]=51761;
squeal_samples[17461]=52837;
squeal_samples[17462]=51968;
squeal_samples[17463]=46679;
squeal_samples[17464]=41516;
squeal_samples[17465]=36693;
squeal_samples[17466]=32175;
squeal_samples[17467]=27943;
squeal_samples[17468]=23991;
squeal_samples[17469]=20287;
squeal_samples[17470]=16825;
squeal_samples[17471]=13578;
squeal_samples[17472]=10551;
squeal_samples[17473]=7709;
squeal_samples[17474]=6174;
squeal_samples[17475]=8865;
squeal_samples[17476]=11826;
squeal_samples[17477]=14669;
squeal_samples[17478]=17382;
squeal_samples[17479]=19980;
squeal_samples[17480]=22465;
squeal_samples[17481]=24832;
squeal_samples[17482]=27107;
squeal_samples[17483]=29272;
squeal_samples[17484]=31345;
squeal_samples[17485]=33326;
squeal_samples[17486]=35221;
squeal_samples[17487]=37026;
squeal_samples[17488]=38753;
squeal_samples[17489]=40403;
squeal_samples[17490]=41974;
squeal_samples[17491]=43489;
squeal_samples[17492]=44914;
squeal_samples[17493]=46295;
squeal_samples[17494]=47603;
squeal_samples[17495]=48856;
squeal_samples[17496]=50056;
squeal_samples[17497]=51196;
squeal_samples[17498]=52293;
squeal_samples[17499]=53126;
squeal_samples[17500]=49373;
squeal_samples[17501]=44040;
squeal_samples[17502]=39055;
squeal_samples[17503]=34383;
squeal_samples[17504]=30011;
squeal_samples[17505]=25924;
squeal_samples[17506]=22099;
squeal_samples[17507]=18516;
squeal_samples[17508]=15166;
squeal_samples[17509]=12028;
squeal_samples[17510]=9100;
squeal_samples[17511]=6398;
squeal_samples[17512]=7319;
squeal_samples[17513]=10349;
squeal_samples[17514]=13245;
squeal_samples[17515]=16035;
squeal_samples[17516]=18680;
squeal_samples[17517]=21231;
squeal_samples[17518]=23650;
squeal_samples[17519]=25972;
squeal_samples[17520]=28190;
squeal_samples[17521]=30308;
squeal_samples[17522]=32336;
squeal_samples[17523]=34270;
squeal_samples[17524]=36119;
squeal_samples[17525]=37888;
squeal_samples[17526]=39577;
squeal_samples[17527]=41188;
squeal_samples[17528]=42729;
squeal_samples[17529]=44201;
squeal_samples[17530]=45600;
squeal_samples[17531]=46942;
squeal_samples[17532]=48224;
squeal_samples[17533]=49450;
squeal_samples[17534]=50620;
squeal_samples[17535]=51740;
squeal_samples[17536]=52810;
squeal_samples[17537]=51945;
squeal_samples[17538]=46655;
squeal_samples[17539]=41490;
squeal_samples[17540]=36669;
squeal_samples[17541]=32151;
squeal_samples[17542]=27917;
squeal_samples[17543]=23970;
squeal_samples[17544]=20259;
squeal_samples[17545]=16803;
squeal_samples[17546]=13552;
squeal_samples[17547]=10527;
squeal_samples[17548]=7686;
squeal_samples[17549]=6148;
squeal_samples[17550]=8841;
squeal_samples[17551]=11803;
squeal_samples[17552]=14641;
squeal_samples[17553]=17362;
squeal_samples[17554]=19952;
squeal_samples[17555]=22443;
squeal_samples[17556]=24806;
squeal_samples[17557]=27084;
squeal_samples[17558]=29245;
squeal_samples[17559]=31323;
squeal_samples[17560]=33301;
squeal_samples[17561]=35194;
squeal_samples[17562]=37006;
squeal_samples[17563]=38723;
squeal_samples[17564]=40384;
squeal_samples[17565]=41947;
squeal_samples[17566]=43462;
squeal_samples[17567]=44895;
squeal_samples[17568]=46264;
squeal_samples[17569]=47584;
squeal_samples[17570]=48828;
squeal_samples[17571]=50031;
squeal_samples[17572]=51174;
squeal_samples[17573]=52265;
squeal_samples[17574]=53261;
squeal_samples[17575]=50161;
squeal_samples[17576]=44778;
squeal_samples[17577]=39740;
squeal_samples[17578]=35023;
squeal_samples[17579]=30609;
squeal_samples[17580]=26482;
squeal_samples[17581]=22616;
squeal_samples[17582]=19003;
squeal_samples[17583]=15617;
squeal_samples[17584]=12453;
squeal_samples[17585]=9489;
squeal_samples[17586]=6719;
squeal_samples[17587]=6961;
squeal_samples[17588]=10009;
squeal_samples[17589]=12919;
squeal_samples[17590]=15713;
squeal_samples[17591]=18377;
squeal_samples[17592]=20932;
squeal_samples[17593]=23372;
squeal_samples[17594]=25703;
squeal_samples[17595]=27933;
squeal_samples[17596]=30058;
squeal_samples[17597]=32100;
squeal_samples[17598]=34038;
squeal_samples[17599]=35904;
squeal_samples[17600]=37677;
squeal_samples[17601]=39373;
squeal_samples[17602]=40997;
squeal_samples[17603]=42538;
squeal_samples[17604]=44022;
squeal_samples[17605]=45426;
squeal_samples[17606]=46779;
squeal_samples[17607]=48066;
squeal_samples[17608]=49297;
squeal_samples[17609]=50469;
squeal_samples[17610]=51596;
squeal_samples[17611]=52668;
squeal_samples[17612]=52858;
squeal_samples[17613]=48105;
squeal_samples[17614]=42854;
squeal_samples[17615]=37935;
squeal_samples[17616]=33337;
squeal_samples[17617]=29030;
squeal_samples[17618]=25000;
squeal_samples[17619]=21233;
squeal_samples[17620]=17702;
squeal_samples[17621]=14400;
squeal_samples[17622]=11315;
squeal_samples[17623]=8424;
squeal_samples[17624]=6124;
squeal_samples[17625]=8113;
squeal_samples[17626]=11110;
squeal_samples[17627]=13978;
squeal_samples[17628]=16721;
squeal_samples[17629]=19344;
squeal_samples[17630]=21851;
squeal_samples[17631]=24246;
squeal_samples[17632]=26543;
squeal_samples[17633]=28733;
squeal_samples[17634]=30832;
squeal_samples[17635]=32829;
squeal_samples[17636]=34746;
squeal_samples[17637]=36567;
squeal_samples[17638]=38317;
squeal_samples[17639]=39976;
squeal_samples[17640]=41576;
squeal_samples[17641]=43094;
squeal_samples[17642]=44549;
squeal_samples[17643]=45932;
squeal_samples[17644]=47260;
squeal_samples[17645]=48520;
squeal_samples[17646]=49738;
squeal_samples[17647]=50884;
squeal_samples[17648]=51994;
squeal_samples[17649]=53048;
squeal_samples[17650]=51503;
squeal_samples[17651]=46083;
squeal_samples[17652]=40962;
squeal_samples[17653]=36162;
squeal_samples[17654]=31682;
squeal_samples[17655]=27472;
squeal_samples[17656]=23552;
squeal_samples[17657]=19873;
squeal_samples[17658]=16429;
squeal_samples[17659]=13211;
squeal_samples[17660]=10198;
squeal_samples[17661]=7379;
squeal_samples[17662]=6346;
squeal_samples[17663]=9238;
squeal_samples[17664]=12188;
squeal_samples[17665]=15011;
squeal_samples[17666]=17705;
squeal_samples[17667]=20290;
squeal_samples[17668]=22755;
squeal_samples[17669]=25109;
squeal_samples[17670]=27364;
squeal_samples[17671]=29523;
squeal_samples[17672]=31574;
squeal_samples[17673]=33550;
squeal_samples[17674]=35422;
squeal_samples[17675]=37223;
squeal_samples[17676]=38935;
squeal_samples[17677]=40575;
squeal_samples[17678]=42138;
squeal_samples[17679]=43633;
squeal_samples[17680]=45067;
squeal_samples[17681]=46423;
squeal_samples[17682]=47730;
squeal_samples[17683]=48973;
squeal_samples[17684]=50161;
squeal_samples[17685]=51301;
squeal_samples[17686]=52382;
squeal_samples[17687]=53212;
squeal_samples[17688]=49452;
squeal_samples[17689]=44111;
squeal_samples[17690]=39110;
squeal_samples[17691]=34440;
squeal_samples[17692]=30055;
squeal_samples[17693]=25963;
squeal_samples[17694]=22127;
squeal_samples[17695]=18545;
squeal_samples[17696]=15183;
squeal_samples[17697]=12048;
squeal_samples[17698]=9103;
squeal_samples[17699]=6407;
squeal_samples[17700]=7320;
squeal_samples[17701]=10354;
squeal_samples[17702]=13245;
squeal_samples[17703]=16024;
squeal_samples[17704]=18679;
squeal_samples[17705]=21214;
squeal_samples[17706]=23641;
squeal_samples[17707]=25952;
squeal_samples[17708]=28173;
squeal_samples[17709]=30291;
squeal_samples[17710]=32312;
squeal_samples[17711]=34255;
squeal_samples[17712]=36092;
squeal_samples[17713]=37864;
squeal_samples[17714]=39544;
squeal_samples[17715]=41163;
squeal_samples[17716]=42693;
squeal_samples[17717]=44168;
squeal_samples[17718]=45566;
squeal_samples[17719]=46906;
squeal_samples[17720]=48192;
squeal_samples[17721]=49410;
squeal_samples[17722]=50581;
squeal_samples[17723]=51699;
squeal_samples[17724]=52770;
squeal_samples[17725]=52476;
squeal_samples[17726]=47399;
squeal_samples[17727]=42183;
squeal_samples[17728]=37310;
squeal_samples[17729]=32744;
squeal_samples[17730]=28479;
squeal_samples[17731]=24480;
squeal_samples[17732]=20746;
squeal_samples[17733]=17241;
squeal_samples[17734]=13969;
squeal_samples[17735]=10907;
squeal_samples[17736]=8046;
squeal_samples[17737]=6076;
squeal_samples[17738]=8457;
squeal_samples[17739]=11439;
squeal_samples[17740]=14288;
squeal_samples[17741]=17020;
squeal_samples[17742]=19630;
squeal_samples[17743]=22122;
squeal_samples[17744]=24510;
squeal_samples[17745]=26787;
squeal_samples[17746]=28964;
squeal_samples[17747]=31049;
squeal_samples[17748]=33039;
squeal_samples[17749]=34939;
squeal_samples[17750]=36758;
squeal_samples[17751]=38493;
squeal_samples[17752]=40149;
squeal_samples[17753]=41733;
squeal_samples[17754]=43243;
squeal_samples[17755]=44685;
squeal_samples[17756]=46066;
squeal_samples[17757]=47383;
squeal_samples[17758]=48645;
squeal_samples[17759]=49844;
squeal_samples[17760]=50993;
squeal_samples[17761]=52091;
squeal_samples[17762]=53143;
squeal_samples[17763]=50821;
squeal_samples[17764]=45387;
squeal_samples[17765]=40308;
squeal_samples[17766]=35549;
squeal_samples[17767]=31102;
squeal_samples[17768]=26933;
squeal_samples[17769]=23041;
squeal_samples[17770]=19392;
squeal_samples[17771]=15979;
squeal_samples[17772]=12790;
squeal_samples[17773]=9797;
squeal_samples[17774]=7008;
squeal_samples[17775]=6561;
squeal_samples[17776]=9584;
squeal_samples[17777]=12511;
squeal_samples[17778]=15314;
squeal_samples[17779]=17999;
squeal_samples[17780]=20563;
squeal_samples[17781]=23021;
squeal_samples[17782]=25357;
squeal_samples[17783]=27603;
squeal_samples[17784]=29742;
squeal_samples[17785]=31798;
squeal_samples[17786]=33747;
squeal_samples[17787]=35618;
squeal_samples[17788]=37401;
squeal_samples[17789]=39111;
squeal_samples[17790]=40739;
squeal_samples[17791]=42297;
squeal_samples[17792]=43777;
squeal_samples[17793]=45202;
squeal_samples[17794]=46557;
squeal_samples[17795]=47849;
squeal_samples[17796]=49090;
squeal_samples[17797]=50271;
squeal_samples[17798]=51401;
squeal_samples[17799]=52481;
squeal_samples[17800]=53040;
squeal_samples[17801]=48726;
squeal_samples[17802]=43432;
squeal_samples[17803]=38473;
squeal_samples[17804]=33837;
squeal_samples[17805]=29487;
squeal_samples[17806]=25431;
squeal_samples[17807]=21632;
squeal_samples[17808]=18071;
squeal_samples[17809]=14743;
squeal_samples[17810]=11626;
squeal_samples[17811]=8719;
squeal_samples[17812]=6169;
squeal_samples[17813]=7675;
squeal_samples[17814]=10684;
squeal_samples[17815]=13563;
squeal_samples[17816]=16325;
squeal_samples[17817]=18961;
squeal_samples[17818]=21487;
squeal_samples[17819]=23900;
squeal_samples[17820]=26194;
squeal_samples[17821]=28414;
squeal_samples[17822]=30509;
squeal_samples[17823]=32529;
squeal_samples[17824]=34448;
squeal_samples[17825]=36287;
squeal_samples[17826]=38042;
squeal_samples[17827]=39717;
squeal_samples[17828]=41318;
squeal_samples[17829]=42849;
squeal_samples[17830]=44309;
squeal_samples[17831]=45704;
squeal_samples[17832]=47034;
squeal_samples[17833]=48311;
squeal_samples[17834]=49526;
squeal_samples[17835]=50692;
squeal_samples[17836]=51798;
squeal_samples[17837]=52865;
squeal_samples[17838]=51995;
squeal_samples[17839]=46686;
squeal_samples[17840]=41525;
squeal_samples[17841]=36684;
squeal_samples[17842]=32161;
squeal_samples[17843]=27927;
squeal_samples[17844]=23965;
squeal_samples[17845]=20259;
squeal_samples[17846]=16786;
squeal_samples[17847]=13541;
squeal_samples[17848]=10502;
squeal_samples[17849]=7663;
squeal_samples[17850]=6113;
squeal_samples[17851]=8804;
squeal_samples[17852]=11764;
squeal_samples[17853]=14600;
squeal_samples[17854]=17316;
squeal_samples[17855]=19912;
squeal_samples[17856]=22392;
squeal_samples[17857]=24760;
squeal_samples[17858]=27027;
squeal_samples[17859]=29194;
squeal_samples[17860]=31266;
squeal_samples[17861]=33244;
squeal_samples[17862]=35134;
squeal_samples[17863]=36946;
squeal_samples[17864]=38660;
squeal_samples[17865]=40316;
squeal_samples[17866]=41885;
squeal_samples[17867]=43392;
squeal_samples[17868]=44828;
squeal_samples[17869]=46197;
squeal_samples[17870]=47510;
squeal_samples[17871]=48761;
squeal_samples[17872]=49954;
squeal_samples[17873]=51099;
squeal_samples[17874]=52189;
squeal_samples[17875]=53185;
squeal_samples[17876]=50082;
squeal_samples[17877]=44694;
squeal_samples[17878]=39662;
squeal_samples[17879]=34939;
squeal_samples[17880]=30526;
squeal_samples[17881]=26398;
squeal_samples[17882]=22531;
squeal_samples[17883]=18915;
squeal_samples[17884]=15533;
squeal_samples[17885]=12365;
squeal_samples[17886]=9404;
squeal_samples[17887]=6631;
squeal_samples[17888]=6869;
squeal_samples[17889]=9919;
squeal_samples[17890]=12830;
squeal_samples[17891]=15624;
squeal_samples[17892]=18288;
squeal_samples[17893]=20846;
squeal_samples[17894]=23282;
squeal_samples[17895]=25607;
squeal_samples[17896]=27846;
squeal_samples[17897]=29963;
squeal_samples[17898]=32007;
squeal_samples[17899]=33950;
squeal_samples[17900]=35808;
squeal_samples[17901]=37583;
squeal_samples[17902]=39280;
squeal_samples[17903]=40898;
squeal_samples[17904]=42450;
squeal_samples[17905]=43926;
squeal_samples[17906]=45338;
squeal_samples[17907]=46684;
squeal_samples[17908]=47969;
squeal_samples[17909]=49207;
squeal_samples[17910]=50373;
squeal_samples[17911]=51509;
squeal_samples[17912]=52570;
squeal_samples[17913]=53134;
squeal_samples[17914]=48803;
squeal_samples[17915]=43509;
squeal_samples[17916]=38536;
squeal_samples[17917]=33899;
squeal_samples[17918]=29544;
squeal_samples[17919]=25480;
squeal_samples[17920]=21672;
squeal_samples[17921]=18110;
squeal_samples[17922]=14775;
squeal_samples[17923]=11659;
squeal_samples[17924]=8738;
squeal_samples[17925]=6190;
squeal_samples[17926]=7690;
squeal_samples[17927]=10696;
squeal_samples[17928]=13578;
squeal_samples[17929]=16334;
squeal_samples[17930]=18971;
squeal_samples[17931]=21492;
squeal_samples[17932]=23905;
squeal_samples[17933]=26206;
squeal_samples[17934]=28408;
squeal_samples[17935]=30512;
squeal_samples[17936]=32520;
squeal_samples[17937]=34446;
squeal_samples[17938]=36278;
squeal_samples[17939]=38031;
squeal_samples[17940]=39708;
squeal_samples[17941]=41309;
squeal_samples[17942]=42838;
squeal_samples[17943]=44302;
squeal_samples[17944]=45686;
squeal_samples[17945]=47027;
squeal_samples[17946]=48294;
squeal_samples[17947]=49512;
squeal_samples[17948]=50671;
squeal_samples[17949]=51777;
squeal_samples[17950]=52844;
squeal_samples[17951]=52544;
squeal_samples[17952]=47455;
squeal_samples[17953]=42237;
squeal_samples[17954]=37353;
squeal_samples[17955]=32783;
squeal_samples[17956]=28500;
squeal_samples[17957]=24502;
squeal_samples[17958]=20758;
squeal_samples[17959]=17256;
squeal_samples[17960]=13975;
squeal_samples[17961]=10907;
squeal_samples[17962]=8037;
squeal_samples[17963]=6068;
squeal_samples[17964]=8444;
squeal_samples[17965]=11425;
squeal_samples[17966]=14268;
squeal_samples[17967]=17000;
squeal_samples[17968]=19605;
squeal_samples[17969]=22103;
squeal_samples[17970]=24477;
squeal_samples[17971]=26759;
squeal_samples[17972]=28934;
squeal_samples[17973]=31017;
squeal_samples[17974]=33008;
squeal_samples[17975]=34899;
squeal_samples[17976]=36723;
squeal_samples[17977]=38447;
squeal_samples[17978]=40112;
squeal_samples[17979]=41686;
squeal_samples[17980]=43202;
squeal_samples[17981]=44640;
squeal_samples[17982]=46018;
squeal_samples[17983]=47340;
squeal_samples[17984]=48591;
squeal_samples[17985]=49794;
squeal_samples[17986]=50946;
squeal_samples[17987]=52037;
squeal_samples[17988]=53095;
squeal_samples[17989]=51531;
squeal_samples[17990]=46106;
squeal_samples[17991]=40975;
squeal_samples[17992]=36169;
squeal_samples[17993]=31677;
squeal_samples[17994]=27470;
squeal_samples[17995]=23536;
squeal_samples[17996]=19852;
squeal_samples[17997]=16402;
squeal_samples[17998]=13175;
squeal_samples[17999]=10162;
squeal_samples[18000]=7337;
squeal_samples[18001]=6303;
squeal_samples[18002]=9192;
squeal_samples[18003]=12137;
squeal_samples[18004]=14950;
squeal_samples[18005]=17654;
squeal_samples[18006]=20232;
squeal_samples[18007]=22695;
squeal_samples[18008]=25048;
squeal_samples[18009]=27299;
squeal_samples[18010]=29454;
squeal_samples[18011]=31511;
squeal_samples[18012]=33477;
squeal_samples[18013]=35350;
squeal_samples[18014]=37152;
squeal_samples[18015]=38858;
squeal_samples[18016]=40497;
squeal_samples[18017]=42062;
squeal_samples[18018]=43552;
squeal_samples[18019]=44980;
squeal_samples[18020]=46344;
squeal_samples[18021]=47647;
squeal_samples[18022]=48888;
squeal_samples[18023]=50078;
squeal_samples[18024]=51206;
squeal_samples[18025]=52298;
squeal_samples[18026]=53279;
squeal_samples[18027]=50175;
squeal_samples[18028]=44778;
squeal_samples[18029]=39728;
squeal_samples[18030]=35008;
squeal_samples[18031]=30582;
squeal_samples[18032]=26449;
squeal_samples[18033]=22580;
squeal_samples[18034]=18953;
squeal_samples[18035]=15565;
squeal_samples[18036]=12390;
squeal_samples[18037]=9430;
squeal_samples[18038]=6643;
squeal_samples[18039]=6890;
squeal_samples[18040]=9925;
squeal_samples[18041]=12838;
squeal_samples[18042]=15628;
squeal_samples[18043]=18290;
squeal_samples[18044]=20844;
squeal_samples[18045]=23282;
squeal_samples[18046]=25610;
squeal_samples[18047]=27834;
squeal_samples[18048]=29966;
squeal_samples[18049]=31995;
squeal_samples[18050]=33942;
squeal_samples[18051]=35798;
squeal_samples[18052]=37568;
squeal_samples[18053]=39269;
squeal_samples[18054]=40877;
squeal_samples[18055]=42431;
squeal_samples[18056]=43903;
squeal_samples[18057]=45317;
squeal_samples[18058]=46661;
squeal_samples[18059]=47950;
squeal_samples[18060]=49176;
squeal_samples[18061]=50350;
squeal_samples[18062]=51477;
squeal_samples[18063]=52548;
squeal_samples[18064]=53102;
squeal_samples[18065]=48782;
squeal_samples[18066]=43470;
squeal_samples[18067]=38509;
squeal_samples[18068]=33861;
squeal_samples[18069]=29516;
squeal_samples[18070]=25440;
squeal_samples[18071]=21639;
squeal_samples[18072]=18074;
squeal_samples[18073]=14735;
squeal_samples[18074]=11622;
squeal_samples[18075]=8700;
squeal_samples[18076]=6151;
squeal_samples[18077]=7648;
squeal_samples[18078]=10658;
squeal_samples[18079]=13539;
squeal_samples[18080]=16291;
squeal_samples[18081]=18933;
squeal_samples[18082]=21449;
squeal_samples[18083]=23862;
squeal_samples[18084]=26161;
squeal_samples[18085]=28367;
squeal_samples[18086]=30466;
squeal_samples[18087]=32480;
squeal_samples[18088]=34400;
squeal_samples[18089]=36235;
squeal_samples[18090]=37989;
squeal_samples[18091]=39663;
squeal_samples[18092]=41267;
squeal_samples[18093]=42789;
squeal_samples[18094]=44252;
squeal_samples[18095]=45645;
squeal_samples[18096]=46976;
squeal_samples[18097]=48251;
squeal_samples[18098]=49465;
squeal_samples[18099]=50624;
squeal_samples[18100]=51739;
squeal_samples[18101]=52790;
squeal_samples[18102]=52500;
squeal_samples[18103]=47403;
squeal_samples[18104]=42189;
squeal_samples[18105]=37305;
squeal_samples[18106]=32733;
squeal_samples[18107]=28460;
squeal_samples[18108]=24449;
squeal_samples[18109]=20712;
squeal_samples[18110]=17205;
squeal_samples[18111]=13929;
squeal_samples[18112]=10856;
squeal_samples[18113]=7990;
squeal_samples[18114]=6017;
squeal_samples[18115]=8404;
squeal_samples[18116]=11372;
squeal_samples[18117]=14230;
squeal_samples[18118]=16950;
squeal_samples[18119]=19563;
squeal_samples[18120]=22050;
squeal_samples[18121]=24430;
squeal_samples[18122]=26710;
squeal_samples[18123]=28884;
squeal_samples[18124]=30971;
squeal_samples[18125]=32955;
squeal_samples[18126]=34856;
squeal_samples[18127]=36668;
squeal_samples[18128]=38403;
squeal_samples[18129]=40061;
squeal_samples[18130]=41636;
squeal_samples[18131]=43156;
squeal_samples[18132]=44594;
squeal_samples[18133]=45972;
squeal_samples[18134]=47287;
squeal_samples[18135]=48546;
squeal_samples[18136]=49748;
squeal_samples[18137]=50899;
squeal_samples[18138]=51988;
squeal_samples[18139]=53045;
squeal_samples[18140]=51484;
squeal_samples[18141]=46056;
squeal_samples[18142]=40927;
squeal_samples[18143]=36119;
squeal_samples[18144]=31630;
squeal_samples[18145]=27420;
squeal_samples[18146]=23489;
squeal_samples[18147]=19802;
squeal_samples[18148]=16352;
squeal_samples[18149]=13127;
squeal_samples[18150]=10114;
squeal_samples[18151]=7288;
squeal_samples[18152]=6255;
squeal_samples[18153]=9141;
squeal_samples[18154]=12094;
squeal_samples[18155]=14903;
squeal_samples[18156]=17604;
squeal_samples[18157]=20183;
squeal_samples[18158]=22647;
squeal_samples[18159]=24999;
squeal_samples[18160]=27250;
squeal_samples[18161]=29405;
squeal_samples[18162]=31463;
squeal_samples[18163]=33426;
squeal_samples[18164]=35304;
squeal_samples[18165]=37103;
squeal_samples[18166]=38806;
squeal_samples[18167]=40453;
squeal_samples[18168]=42008;
squeal_samples[18169]=43506;
squeal_samples[18170]=44932;
squeal_samples[18171]=46293;
squeal_samples[18172]=47600;
squeal_samples[18173]=48838;
squeal_samples[18174]=50029;
squeal_samples[18175]=51159;
squeal_samples[18176]=52247;
squeal_samples[18177]=53232;
squeal_samples[18178]=50125;
squeal_samples[18179]=44729;
squeal_samples[18180]=39681;
squeal_samples[18181]=34957;
squeal_samples[18182]=30536;
squeal_samples[18183]=26396;
squeal_samples[18184]=22535;
squeal_samples[18185]=18902;
squeal_samples[18186]=15517;
squeal_samples[18187]=12343;
squeal_samples[18188]=9376;
squeal_samples[18189]=6600;
squeal_samples[18190]=6837;
squeal_samples[18191]=9879;
squeal_samples[18192]=12788;
squeal_samples[18193]=15579;
squeal_samples[18194]=18241;
squeal_samples[18195]=20796;
squeal_samples[18196]=23233;
squeal_samples[18197]=25560;
squeal_samples[18198]=27788;
squeal_samples[18199]=29912;
squeal_samples[18200]=31951;
squeal_samples[18201]=33891;
squeal_samples[18202]=35749;
squeal_samples[18203]=37521;
squeal_samples[18204]=39217;
squeal_samples[18205]=40831;
squeal_samples[18206]=42381;
squeal_samples[18207]=43854;
squeal_samples[18208]=45269;
squeal_samples[18209]=46612;
squeal_samples[18210]=47900;
squeal_samples[18211]=49128;
squeal_samples[18212]=50301;
squeal_samples[18213]=51428;
squeal_samples[18214]=52500;
squeal_samples[18215]=53052;
squeal_samples[18216]=48732;
squeal_samples[18217]=43423;
squeal_samples[18218]=38459;
squeal_samples[18219]=33814;
squeal_samples[18220]=29464;
squeal_samples[18221]=25393;
squeal_samples[18222]=21590;
squeal_samples[18223]=18024;
squeal_samples[18224]=14689;
squeal_samples[18225]=11568;
squeal_samples[18226]=8656;
squeal_samples[18227]=6099;
squeal_samples[18228]=7600;
squeal_samples[18229]=10609;
squeal_samples[18230]=13489;
squeal_samples[18231]=16245;
squeal_samples[18232]=18880;
squeal_samples[18233]=21403;
squeal_samples[18234]=23811;
squeal_samples[18235]=26113;
squeal_samples[18236]=28319;
squeal_samples[18237]=30415;
squeal_samples[18238]=32433;
squeal_samples[18239]=34349;
squeal_samples[18240]=36188;
squeal_samples[18241]=37938;
squeal_samples[18242]=39616;
squeal_samples[18243]=41217;
squeal_samples[18244]=42739;
squeal_samples[18245]=44204;
squeal_samples[18246]=45595;
squeal_samples[18247]=46928;
squeal_samples[18248]=48201;
squeal_samples[18249]=49415;
squeal_samples[18250]=50576;
squeal_samples[18251]=51687;
squeal_samples[18252]=52744;
squeal_samples[18253]=52919;
squeal_samples[18254]=48150;
squeal_samples[18255]=42883;
squeal_samples[18256]=37952;
squeal_samples[18257]=33334;
squeal_samples[18258]=29020;
squeal_samples[18259]=24969;
squeal_samples[18260]=21201;
squeal_samples[18261]=17657;
squeal_samples[18262]=14344;
squeal_samples[18263]=11250;
squeal_samples[18264]=8345;
squeal_samples[18265]=6042;
squeal_samples[18266]=8019;
squeal_samples[18267]=11012;
squeal_samples[18268]=13872;
squeal_samples[18269]=16617;
squeal_samples[18270]=19235;
squeal_samples[18271]=21739;
squeal_samples[18272]=24134;
squeal_samples[18273]=26418;
squeal_samples[18274]=28611;
squeal_samples[18275]=30696;
squeal_samples[18276]=32697;
squeal_samples[18277]=34604;
squeal_samples[18278]=36428;
squeal_samples[18279]=38173;
squeal_samples[18280]=39834;
squeal_samples[18281]=41428;
squeal_samples[18282]=42940;
squeal_samples[18283]=44395;
squeal_samples[18284]=45781;
squeal_samples[18285]=47097;
squeal_samples[18286]=48366;
squeal_samples[18287]=49568;
squeal_samples[18288]=50724;
squeal_samples[18289]=51825;
squeal_samples[18290]=52879;
squeal_samples[18291]=52577;
squeal_samples[18292]=47479;
squeal_samples[18293]=42252;
squeal_samples[18294]=37357;
squeal_samples[18295]=32781;
squeal_samples[18296]=28493;
squeal_samples[18297]=24490;
squeal_samples[18298]=20738;
squeal_samples[18299]=17230;
squeal_samples[18300]=13939;
squeal_samples[18301]=10874;
squeal_samples[18302]=7995;
squeal_samples[18303]=6025;
squeal_samples[18304]=8398;
squeal_samples[18305]=11375;
squeal_samples[18306]=14218;
squeal_samples[18307]=16942;
squeal_samples[18308]=19546;
squeal_samples[18309]=22041;
squeal_samples[18310]=24415;
squeal_samples[18311]=26693;
squeal_samples[18312]=28866;
squeal_samples[18313]=30947;
squeal_samples[18314]=32932;
squeal_samples[18315]=34833;
squeal_samples[18316]=36643;
squeal_samples[18317]=38377;
squeal_samples[18318]=40028;
squeal_samples[18319]=41612;
squeal_samples[18320]=43117;
squeal_samples[18321]=44563;
squeal_samples[18322]=45936;
squeal_samples[18323]=47253;
squeal_samples[18324]=48511;
squeal_samples[18325]=49708;
squeal_samples[18326]=50859;
squeal_samples[18327]=51949;
squeal_samples[18328]=53003;
squeal_samples[18329]=52118;
squeal_samples[18330]=46794;
squeal_samples[18331]=41607;
squeal_samples[18332]=36762;
squeal_samples[18333]=32217;
squeal_samples[18334]=27968;
squeal_samples[18335]=23991;
squeal_samples[18336]=20278;
squeal_samples[18337]=16791;
squeal_samples[18338]=13538;
squeal_samples[18339]=10491;
squeal_samples[18340]=7636;
squeal_samples[18341]=6087;
squeal_samples[18342]=8768;
squeal_samples[18343]=11725;
squeal_samples[18344]=14555;
squeal_samples[18345]=17266;
squeal_samples[18346]=19853;
squeal_samples[18347]=22334;
squeal_samples[18348]=24689;
squeal_samples[18349]=26958;
squeal_samples[18350]=29120;
squeal_samples[18351]=31190;
squeal_samples[18352]=33163;
squeal_samples[18353]=35054;
squeal_samples[18354]=36853;
squeal_samples[18355]=38576;
squeal_samples[18356]=40218;
squeal_samples[18357]=41794;
squeal_samples[18358]=43289;
squeal_samples[18359]=44725;
squeal_samples[18360]=46091;
squeal_samples[18361]=47399;
squeal_samples[18362]=48651;
squeal_samples[18363]=49843;
squeal_samples[18364]=50987;
squeal_samples[18365]=52074;
squeal_samples[18366]=53114;
squeal_samples[18367]=51554;
squeal_samples[18368]=46117;
squeal_samples[18369]=40972;
squeal_samples[18370]=36167;
squeal_samples[18371]=31657;
squeal_samples[18372]=27445;
squeal_samples[18373]=23505;
squeal_samples[18374]=19817;
squeal_samples[18375]=16359;
squeal_samples[18376]=13137;
squeal_samples[18377]=10106;
squeal_samples[18378]=7284;
squeal_samples[18379]=6236;
squeal_samples[18380]=9133;
squeal_samples[18381]=12068;
squeal_samples[18382]=14894;
squeal_samples[18383]=17580;
squeal_samples[18384]=20163;
squeal_samples[18385]=22618;
squeal_samples[18386]=24977;
squeal_samples[18387]=27217;
squeal_samples[18388]=29377;
squeal_samples[18389]=31425;
squeal_samples[18390]=33392;
squeal_samples[18391]=35268;
squeal_samples[18392]=37059;
squeal_samples[18393]=38775;
squeal_samples[18394]=40405;
squeal_samples[18395]=41974;
squeal_samples[18396]=43460;
squeal_samples[18397]=44886;
squeal_samples[18398]=46248;
squeal_samples[18399]=47549;
squeal_samples[18400]=48791;
squeal_samples[18401]=49977;
squeal_samples[18402]=51110;
squeal_samples[18403]=52192;
squeal_samples[18404]=53230;
squeal_samples[18405]=50888;
squeal_samples[18406]=45441;
squeal_samples[18407]=40342;
squeal_samples[18408]=35570;
squeal_samples[18409]=31111;
squeal_samples[18410]=26925;
squeal_samples[18411]=23018;
squeal_samples[18412]=19357;
squeal_samples[18413]=15935;
squeal_samples[18414]=12732;
squeal_samples[18415]=9731;
squeal_samples[18416]=6934;
squeal_samples[18417]=6480;
squeal_samples[18418]=9495;
squeal_samples[18419]=12416;
squeal_samples[18420]=15221;
squeal_samples[18421]=17898;
squeal_samples[18422]=20460;
squeal_samples[18423]=22909;
squeal_samples[18424]=25244;
squeal_samples[18425]=27483;
squeal_samples[18426]=29625;
squeal_samples[18427]=31662;
squeal_samples[18428]=33619;
squeal_samples[18429]=35482;
squeal_samples[18430]=37267;
squeal_samples[18431]=38964;
squeal_samples[18432]=40599;
squeal_samples[18433]=42147;
squeal_samples[18434]=43629;
squeal_samples[18435]=45049;
squeal_samples[18436]=46400;
squeal_samples[18437]=47698;
squeal_samples[18438]=48928;
squeal_samples[18439]=50108;
squeal_samples[18440]=51234;
squeal_samples[18441]=52310;
squeal_samples[18442]=53292;
squeal_samples[18443]=50177;
squeal_samples[18444]=44771;
squeal_samples[18445]=39715;
squeal_samples[18446]=34985;
squeal_samples[18447]=30557;
squeal_samples[18448]=26411;
squeal_samples[18449]=22537;
squeal_samples[18450]=18905;
squeal_samples[18451]=15511;
squeal_samples[18452]=12333;
squeal_samples[18453]=9362;
squeal_samples[18454]=6581;
squeal_samples[18455]=6820;
squeal_samples[18456]=9847;
squeal_samples[18457]=12768;
squeal_samples[18458]=15547;
squeal_samples[18459]=18212;
squeal_samples[18460]=20759;
squeal_samples[18461]=23192;
squeal_samples[18462]=25522;
squeal_samples[18463]=27741;
squeal_samples[18464]=29873;
squeal_samples[18465]=31900;
squeal_samples[18466]=33844;
squeal_samples[18467]=35700;
squeal_samples[18468]=37468;
squeal_samples[18469]=39163;
squeal_samples[18470]=40777;
squeal_samples[18471]=42329;
squeal_samples[18472]=43798;
squeal_samples[18473]=45211;
squeal_samples[18474]=46553;
squeal_samples[18475]=47840;
squeal_samples[18476]=49070;
squeal_samples[18477]=50242;
squeal_samples[18478]=51360;
squeal_samples[18479]=52438;
squeal_samples[18480]=53246;
squeal_samples[18481]=49469;
squeal_samples[18482]=44106;
squeal_samples[18483]=39095;
squeal_samples[18484]=34401;
squeal_samples[18485]=30009;
squeal_samples[18486]=25898;
squeal_samples[18487]=22058;
squeal_samples[18488]=18459;
squeal_samples[18489]=15089;
squeal_samples[18490]=11944;
squeal_samples[18491]=8987;
squeal_samples[18492]=6280;
squeal_samples[18493]=7188;
squeal_samples[18494]=10216;
squeal_samples[18495]=13103;
squeal_samples[18496]=15875;
squeal_samples[18497]=18524;
squeal_samples[18498]=21062;
squeal_samples[18499]=23479;
squeal_samples[18500]=25791;
squeal_samples[18501]=28000;
squeal_samples[18502]=30122;
squeal_samples[18503]=32137;
squeal_samples[18504]=34071;
squeal_samples[18505]=35914;
squeal_samples[18506]=37675;
squeal_samples[18507]=39355;
squeal_samples[18508]=40969;
squeal_samples[18509]=42496;
squeal_samples[18510]=43970;
squeal_samples[18511]=45368;
squeal_samples[18512]=46705;
squeal_samples[18513]=47987;
squeal_samples[18514]=49202;
squeal_samples[18515]=50372;
squeal_samples[18516]=51485;
squeal_samples[18517]=52554;
squeal_samples[18518]=53095;
squeal_samples[18519]=48769;
squeal_samples[18520]=43455;
squeal_samples[18521]=38478;
squeal_samples[18522]=33827;
squeal_samples[18523]=29466;
squeal_samples[18524]=25395;
squeal_samples[18525]=21575;
squeal_samples[18526]=18015;
squeal_samples[18527]=14668;
squeal_samples[18528]=11552;
squeal_samples[18529]=8621;
squeal_samples[18530]=6071;
squeal_samples[18531]=7564;
squeal_samples[18532]=10570;
squeal_samples[18533]=13447;
squeal_samples[18534]=16197;
squeal_samples[18535]=18834;
squeal_samples[18536]=21351;
squeal_samples[18537]=23764;
squeal_samples[18538]=26055;
squeal_samples[18539]=28265;
squeal_samples[18540]=30360;
squeal_samples[18541]=32371;
squeal_samples[18542]=34292;
squeal_samples[18543]=36123;
squeal_samples[18544]=37881;
squeal_samples[18545]=39547;
squeal_samples[18546]=41152;
squeal_samples[18547]=42675;
squeal_samples[18548]=44134;
squeal_samples[18549]=45527;
squeal_samples[18550]=46853;
squeal_samples[18551]=48127;
squeal_samples[18552]=49342;
squeal_samples[18553]=50500;
squeal_samples[18554]=51609;
squeal_samples[18555]=52665;
squeal_samples[18556]=53209;
squeal_samples[18557]=48869;
squeal_samples[18558]=43553;
squeal_samples[18559]=38567;
squeal_samples[18560]=33912;
squeal_samples[18561]=29542;
squeal_samples[18562]=25461;
squeal_samples[18563]=21648;
squeal_samples[18564]=18069;
squeal_samples[18565]=14729;
squeal_samples[18566]=11597;
squeal_samples[18567]=8670;
squeal_samples[18568]=6112;
squeal_samples[18569]=7599;
squeal_samples[18570]=10610;
squeal_samples[18571]=13479;
squeal_samples[18572]=16237;
squeal_samples[18573]=18869;
squeal_samples[18574]=21381;
squeal_samples[18575]=23791;
squeal_samples[18576]=26080;
squeal_samples[18577]=28290;
squeal_samples[18578]=30387;
squeal_samples[18579]=32395;
squeal_samples[18580]=34313;
squeal_samples[18581]=36144;
squeal_samples[18582]=37893;
squeal_samples[18583]=39565;
squeal_samples[18584]=41163;
squeal_samples[18585]=42694;
squeal_samples[18586]=44141;
squeal_samples[18587]=45541;
squeal_samples[18588]=46865;
squeal_samples[18589]=48133;
squeal_samples[18590]=49349;
squeal_samples[18591]=50506;
squeal_samples[18592]=51616;
squeal_samples[18593]=52673;
squeal_samples[18594]=53212;
squeal_samples[18595]=48876;
squeal_samples[18596]=43545;
squeal_samples[18597]=38579;
squeal_samples[18598]=33904;
squeal_samples[18599]=29550;
squeal_samples[18600]=25463;
squeal_samples[18601]=21645;
squeal_samples[18602]=18071;
squeal_samples[18603]=14719;
squeal_samples[18604]=11598;
squeal_samples[18605]=8660;
squeal_samples[18606]=6113;
squeal_samples[18607]=7597;
squeal_samples[18608]=10601;
squeal_samples[18609]=13475;
squeal_samples[18610]=16228;
squeal_samples[18611]=18862;
squeal_samples[18612]=21377;
squeal_samples[18613]=23779;
squeal_samples[18614]=26078;
squeal_samples[18615]=28280;
squeal_samples[18616]=30381;
squeal_samples[18617]=32383;
squeal_samples[18618]=34305;
squeal_samples[18619]=36132;
squeal_samples[18620]=37887;
squeal_samples[18621]=39556;
squeal_samples[18622]=41154;
squeal_samples[18623]=42677;
squeal_samples[18624]=44138;
squeal_samples[18625]=45527;
squeal_samples[18626]=46857;
squeal_samples[18627]=48129;
squeal_samples[18628]=49338;
squeal_samples[18629]=50498;
squeal_samples[18630]=51606;
squeal_samples[18631]=52661;
squeal_samples[18632]=53202;
squeal_samples[18633]=48859;
squeal_samples[18634]=43545;
squeal_samples[18635]=38560;
squeal_samples[18636]=33895;
squeal_samples[18637]=29538;
squeal_samples[18638]=25448;
squeal_samples[18639]=21638;
squeal_samples[18640]=18057;
squeal_samples[18641]=14720;
squeal_samples[18642]=11577;
squeal_samples[18643]=8662;
squeal_samples[18644]=6094;
squeal_samples[18645]=7588;
squeal_samples[18646]=10588;
squeal_samples[18647]=13468;
squeal_samples[18648]=16214;
squeal_samples[18649]=18854;
squeal_samples[18650]=21364;
squeal_samples[18651]=23772;
squeal_samples[18652]=26068;
squeal_samples[18653]=28269;
squeal_samples[18654]=30369;
squeal_samples[18655]=32375;
squeal_samples[18656]=34293;
squeal_samples[18657]=36126;
squeal_samples[18658]=37873;
squeal_samples[18659]=39546;
squeal_samples[18660]=41139;
squeal_samples[18661]=42666;
squeal_samples[18662]=44126;
squeal_samples[18663]=45513;
squeal_samples[18664]=46848;
squeal_samples[18665]=48112;
squeal_samples[18666]=49330;
squeal_samples[18667]=50482;
squeal_samples[18668]=51596;
squeal_samples[18669]=52649;
squeal_samples[18670]=53188;
squeal_samples[18671]=48848;
squeal_samples[18672]=43532;
squeal_samples[18673]=38547;
squeal_samples[18674]=33891;
squeal_samples[18675]=29521;
squeal_samples[18676]=25440;
squeal_samples[18677]=21622;
squeal_samples[18678]=18048;
squeal_samples[18679]=14705;
squeal_samples[18680]=11567;
squeal_samples[18681]=8646;
squeal_samples[18682]=6085;
squeal_samples[18683]=7574;
squeal_samples[18684]=10578;
squeal_samples[18685]=13452;
squeal_samples[18686]=16207;
squeal_samples[18687]=18835;
squeal_samples[18688]=21358;
squeal_samples[18689]=23756;
squeal_samples[18690]=26057;
squeal_samples[18691]=28256;
squeal_samples[18692]=30357;
squeal_samples[18693]=32363;
squeal_samples[18694]=34280;
squeal_samples[18695]=36114;
squeal_samples[18696]=37861;
squeal_samples[18697]=39532;
squeal_samples[18698]=41130;
squeal_samples[18699]=42650;
squeal_samples[18700]=44116;
squeal_samples[18701]=45500;
squeal_samples[18702]=46834;
squeal_samples[18703]=48103;
squeal_samples[18704]=49314;
squeal_samples[18705]=50473;
squeal_samples[18706]=51580;
squeal_samples[18707]=52640;
squeal_samples[18708]=53172;
squeal_samples[18709]=48839;
squeal_samples[18710]=43518;
squeal_samples[18711]=38536;
squeal_samples[18712]=33876;
squeal_samples[18713]=29512;
squeal_samples[18714]=25424;
squeal_samples[18715]=21613;
squeal_samples[18716]=18035;
squeal_samples[18717]=14690;
squeal_samples[18718]=11559;
squeal_samples[18719]=8631;
squeal_samples[18720]=6074;
squeal_samples[18721]=7560;
squeal_samples[18722]=10566;
squeal_samples[18723]=13441;
squeal_samples[18724]=16194;
squeal_samples[18725]=18822;
squeal_samples[18726]=21347;
squeal_samples[18727]=23741;
squeal_samples[18728]=26048;
squeal_samples[18729]=28242;
squeal_samples[18730]=30344;
squeal_samples[18731]=32352;
squeal_samples[18732]=34266;
squeal_samples[18733]=36104;
squeal_samples[18734]=37847;
squeal_samples[18735]=39522;
squeal_samples[18736]=41114;
squeal_samples[18737]=42642;
squeal_samples[18738]=44100;
squeal_samples[18739]=45491;
squeal_samples[18740]=46821;
squeal_samples[18741]=48089;
squeal_samples[18742]=49305;
squeal_samples[18743]=50456;
squeal_samples[18744]=51573;
squeal_samples[18745]=52624;
squeal_samples[18746]=53162;
squeal_samples[18747]=48827;
squeal_samples[18748]=43502;
squeal_samples[18749]=38527;
squeal_samples[18750]=33863;
squeal_samples[18751]=29499;
squeal_samples[18752]=25414;
squeal_samples[18753]=21598;
squeal_samples[18754]=18023;
squeal_samples[18755]=14679;
squeal_samples[18756]=11545;
squeal_samples[18757]=8620;
squeal_samples[18758]=6061;
squeal_samples[18759]=7549;
squeal_samples[18760]=10552;
squeal_samples[18761]=13430;
squeal_samples[18762]=16179;
squeal_samples[18763]=18814;
squeal_samples[18764]=21330;
squeal_samples[18765]=23734;
squeal_samples[18766]=26031;
squeal_samples[18767]=28232;
squeal_samples[18768]=30332;
squeal_samples[18769]=32338;
squeal_samples[18770]=34256;
squeal_samples[18771]=36089;
squeal_samples[18772]=37838;
squeal_samples[18773]=39506;
squeal_samples[18774]=41105;
squeal_samples[18775]=42627;
squeal_samples[18776]=44089;
squeal_samples[18777]=45479;
squeal_samples[18778]=46807;
squeal_samples[18779]=48078;
squeal_samples[18780]=49292;
squeal_samples[18781]=50446;
squeal_samples[18782]=51557;
squeal_samples[18783]=52615;
squeal_samples[18784]=53147;
squeal_samples[18785]=48816;
squeal_samples[18786]=43491;
squeal_samples[18787]=38512;
squeal_samples[18788]=33854;
squeal_samples[18789]=29483;
squeal_samples[18790]=25405;
squeal_samples[18791]=21584;
squeal_samples[18792]=18010;
squeal_samples[18793]=14670;
squeal_samples[18794]=11528;
squeal_samples[18795]=8612;
squeal_samples[18796]=6045;
squeal_samples[18797]=7540;
squeal_samples[18798]=10537;
squeal_samples[18799]=13420;
squeal_samples[18800]=16166;
squeal_samples[18801]=18800;
squeal_samples[18802]=21321;
squeal_samples[18803]=23718;
squeal_samples[18804]=26021;
squeal_samples[18805]=28220;
squeal_samples[18806]=30317;
squeal_samples[18807]=32329;
squeal_samples[18808]=34242;
squeal_samples[18809]=36077;
squeal_samples[18810]=37825;
squeal_samples[18811]=39495;
squeal_samples[18812]=41092;
squeal_samples[18813]=42616;
squeal_samples[18814]=44075;
squeal_samples[18815]=45468;
squeal_samples[18816]=46793;
squeal_samples[18817]=48070;
squeal_samples[18818]=49273;
squeal_samples[18819]=50440;
squeal_samples[18820]=51541;
squeal_samples[18821]=52603;
squeal_samples[18822]=53137;
squeal_samples[18823]=48799;
squeal_samples[18824]=43484;
squeal_samples[18825]=38497;
squeal_samples[18826]=33842;
squeal_samples[18827]=29472;
squeal_samples[18828]=25390;
squeal_samples[18829]=21574;
squeal_samples[18830]=17998;
squeal_samples[18831]=14656;
squeal_samples[18832]=11518;
squeal_samples[18833]=8598;
squeal_samples[18834]=6034;
squeal_samples[18835]=7526;
squeal_samples[18836]=10526;
squeal_samples[18837]=13407;
squeal_samples[18838]=16153;
squeal_samples[18839]=18790;
squeal_samples[18840]=21307;
squeal_samples[18841]=23706;
squeal_samples[18842]=26009;
squeal_samples[18843]=28206;
squeal_samples[18844]=30307;
squeal_samples[18845]=32316;
squeal_samples[18846]=34230;
squeal_samples[18847]=36063;
squeal_samples[18848]=37815;
squeal_samples[18849]=39480;
squeal_samples[18850]=41082;
squeal_samples[18851]=42602;
squeal_samples[18852]=44064;
squeal_samples[18853]=45455;
squeal_samples[18854]=46781;
squeal_samples[18855]=48057;
squeal_samples[18856]=49262;
squeal_samples[18857]=50426;
squeal_samples[18858]=51530;
squeal_samples[18859]=52591;
squeal_samples[18860]=53123;
squeal_samples[18861]=48791;
squeal_samples[18862]=43465;
squeal_samples[18863]=38490;
squeal_samples[18864]=33826;
squeal_samples[18865]=29462;
squeal_samples[18866]=25378;
squeal_samples[18867]=21559;
squeal_samples[18868]=17989;
squeal_samples[18869]=14640;
squeal_samples[18870]=11509;
squeal_samples[18871]=8583;
squeal_samples[18872]=6023;
squeal_samples[18873]=7514;
squeal_samples[18874]=10514;
squeal_samples[18875]=13393;
squeal_samples[18876]=16143;
squeal_samples[18877]=18775;
squeal_samples[18878]=21297;
squeal_samples[18879]=23692;
squeal_samples[18880]=25999;
squeal_samples[18881]=28190;
squeal_samples[18882]=30300;
squeal_samples[18883]=32297;
squeal_samples[18884]=34223;
squeal_samples[18885]=36048;
squeal_samples[18886]=37802;
squeal_samples[18887]=39471;
squeal_samples[18888]=41065;
squeal_samples[18889]=42593;
squeal_samples[18890]=44050;
squeal_samples[18891]=45441;
squeal_samples[18892]=46773;
squeal_samples[18893]=48038;
squeal_samples[18894]=49257;
squeal_samples[18895]=50406;
squeal_samples[18896]=51523;
squeal_samples[18897]=52574;
squeal_samples[18898]=53378;
squeal_samples[18899]=49588;
squeal_samples[18900]=44209;
squeal_samples[18901]=39182;
squeal_samples[18902]=34471;
squeal_samples[18903]=30069;
squeal_samples[18904]=25945;
squeal_samples[18905]=22093;
squeal_samples[18906]=18478;
squeal_samples[18907]=15102;
squeal_samples[18908]=11942;
squeal_samples[18909]=8982;
squeal_samples[18910]=6269;
squeal_samples[18911]=7166;
squeal_samples[18912]=10189;
squeal_samples[18913]=13075;
squeal_samples[18914]=15844;
squeal_samples[18915]=18485;
squeal_samples[18916]=21017;
squeal_samples[18917]=23432;
squeal_samples[18918]=25740;
squeal_samples[18919]=27948;
squeal_samples[18920]=30060;
squeal_samples[18921]=32078;
squeal_samples[18922]=34006;
squeal_samples[18923]=35842;
squeal_samples[18924]=37606;
squeal_samples[18925]=39282;
squeal_samples[18926]=40888;
squeal_samples[18927]=42421;
squeal_samples[18928]=43886;
squeal_samples[18929]=45284;
squeal_samples[18930]=46615;
squeal_samples[18931]=47896;
squeal_samples[18932]=49107;
squeal_samples[18933]=50282;
squeal_samples[18934]=51383;
squeal_samples[18935]=52459;
squeal_samples[18936]=53410;
squeal_samples[18937]=50289;
squeal_samples[18938]=44865;
squeal_samples[18939]=39793;
squeal_samples[18940]=35048;
squeal_samples[18941]=30602;
squeal_samples[18942]=26446;
squeal_samples[18943]=22555;
squeal_samples[18944]=18920;
squeal_samples[18945]=15505;
squeal_samples[18946]=12322;
squeal_samples[18947]=9340;
squeal_samples[18948]=6554;
squeal_samples[18949]=6776;
squeal_samples[18950]=9808;
squeal_samples[18951]=12720;
squeal_samples[18952]=15489;
squeal_samples[18953]=18159;
squeal_samples[18954]=20696;
squeal_samples[18955]=23129;
squeal_samples[18956]=25450;
squeal_samples[18957]=27669;
squeal_samples[18958]=29794;
squeal_samples[18959]=31821;
squeal_samples[18960]=33759;
squeal_samples[18961]=35610;
squeal_samples[18962]=37379;
squeal_samples[18963]=39066;
squeal_samples[18964]=40684;
squeal_samples[18965]=42224;
squeal_samples[18966]=43696;
squeal_samples[18967]=45102;
squeal_samples[18968]=46446;
squeal_samples[18969]=47731;
squeal_samples[18970]=48955;
squeal_samples[18971]=50126;
squeal_samples[18972]=51243;
squeal_samples[18973]=52312;
squeal_samples[18974]=53337;
squeal_samples[18975]=50979;
squeal_samples[18976]=45514;
squeal_samples[18977]=40397;
squeal_samples[18978]=35612;
squeal_samples[18979]=31128;
squeal_samples[18980]=26938;
squeal_samples[18981]=23017;
squeal_samples[18982]=19344;
squeal_samples[18983]=15915;
squeal_samples[18984]=12697;
squeal_samples[18985]=9689;
squeal_samples[18986]=6878;
squeal_samples[18987]=6420;
squeal_samples[18988]=9429;
squeal_samples[18989]=12345;
squeal_samples[18990]=15145;
squeal_samples[18991]=17815;
squeal_samples[18992]=20374;
squeal_samples[18993]=22821;
squeal_samples[18994]=25150;
squeal_samples[18995]=27387;
squeal_samples[18996]=29519;
squeal_samples[18997]=31561;
squeal_samples[18998]=33507;
squeal_samples[18999]=35376;
squeal_samples[19000]=37149;
squeal_samples[19001]=38849;
squeal_samples[19002]=40469;
squeal_samples[19003]=42024;
squeal_samples[19004]=43503;
squeal_samples[19005]=44923;
squeal_samples[19006]=46265;
squeal_samples[19007]=47561;
squeal_samples[19008]=48791;
squeal_samples[19009]=49971;
squeal_samples[19010]=51098;
squeal_samples[19011]=52166;
squeal_samples[19012]=53201;
squeal_samples[19013]=51619;
squeal_samples[19014]=46161;
squeal_samples[19015]=41010;
squeal_samples[19016]=36181;
squeal_samples[19017]=31667;
squeal_samples[19018]=27436;
squeal_samples[19019]=23481;
squeal_samples[19020]=19779;
squeal_samples[19021]=16314;
squeal_samples[19022]=13078;
squeal_samples[19023]=10044;
squeal_samples[19024]=7210;
squeal_samples[19025]=6157;
squeal_samples[19026]=9040;
squeal_samples[19027]=11978;
squeal_samples[19028]=14787;
squeal_samples[19029]=17479;
squeal_samples[19030]=20051;
squeal_samples[19031]=22510;
squeal_samples[19032]=24857;
squeal_samples[19033]=27102;
squeal_samples[19034]=29247;
squeal_samples[19035]=31298;
squeal_samples[19036]=33257;
squeal_samples[19037]=35130;
squeal_samples[19038]=36919;
squeal_samples[19039]=38631;
squeal_samples[19040]=40262;
squeal_samples[19041]=41821;
squeal_samples[19042]=43313;
squeal_samples[19043]=44734;
squeal_samples[19044]=46093;
squeal_samples[19045]=47389;
squeal_samples[19046]=48628;
squeal_samples[19047]=49814;
squeal_samples[19048]=50939;
squeal_samples[19049]=52030;
squeal_samples[19050]=53056;
squeal_samples[19051]=52166;
squeal_samples[19052]=46817;
squeal_samples[19053]=41620;
squeal_samples[19054]=36753;
squeal_samples[19055]=32201;
squeal_samples[19056]=27939;
squeal_samples[19057]=23948;
squeal_samples[19058]=20217;
squeal_samples[19059]=16726;
squeal_samples[19060]=13455;
squeal_samples[19061]=10397;
squeal_samples[19062]=7540;
squeal_samples[19063]=5975;
squeal_samples[19064]=8655;
squeal_samples[19065]=11604;
squeal_samples[19066]=14430;
squeal_samples[19067]=17134;
squeal_samples[19068]=19725;
squeal_samples[19069]=22192;
squeal_samples[19070]=24560;
squeal_samples[19071]=26809;
squeal_samples[19072]=28980;
squeal_samples[19073]=31030;
squeal_samples[19074]=33011;
squeal_samples[19075]=34887;
squeal_samples[19076]=36691;
squeal_samples[19077]=38407;
squeal_samples[19078]=40049;
squeal_samples[19079]=41619;
squeal_samples[19080]=43115;
squeal_samples[19081]=44550;
squeal_samples[19082]=45911;
squeal_samples[19083]=47220;
squeal_samples[19084]=48465;
squeal_samples[19085]=49651;
squeal_samples[19086]=50796;
squeal_samples[19087]=51882;
squeal_samples[19088]=52917;
squeal_samples[19089]=52603;
squeal_samples[19090]=47483;
squeal_samples[19091]=42246;
squeal_samples[19092]=37330;
squeal_samples[19093]=32739;
squeal_samples[19094]=28442;
squeal_samples[19095]=24420;
squeal_samples[19096]=20660;
squeal_samples[19097]=17138;
squeal_samples[19098]=13839;
squeal_samples[19099]=10760;
squeal_samples[19100]=7875;
squeal_samples[19101]=5889;
squeal_samples[19102]=8260;
squeal_samples[19103]=11235;
squeal_samples[19104]=14073;
squeal_samples[19105]=16794;
squeal_samples[19106]=19388;
squeal_samples[19107]=21882;
squeal_samples[19108]=24247;
squeal_samples[19109]=26528;
squeal_samples[19110]=28694;
squeal_samples[19111]=30769;
squeal_samples[19112]=32756;
squeal_samples[19113]=34649;
squeal_samples[19114]=36456;
squeal_samples[19115]=38188;
squeal_samples[19116]=39836;
squeal_samples[19117]=41416;
squeal_samples[19118]=42921;
squeal_samples[19119]=44356;
squeal_samples[19120]=45732;
squeal_samples[19121]=47045;
squeal_samples[19122]=48298;
squeal_samples[19123]=49501;
squeal_samples[19124]=50641;
squeal_samples[19125]=51733;
squeal_samples[19126]=52782;
squeal_samples[19127]=52940;
squeal_samples[19128]=48154;
squeal_samples[19129]=42866;
squeal_samples[19130]=37918;
squeal_samples[19131]=33285;
squeal_samples[19132]=28953;
squeal_samples[19133]=24893;
squeal_samples[19134]=21108;
squeal_samples[19135]=17550;
squeal_samples[19136]=14234;
squeal_samples[19137]=11115;
squeal_samples[19138]=8210;
squeal_samples[19139]=5894;
squeal_samples[19140]=7867;
squeal_samples[19141]=10858;
squeal_samples[19142]=13710;
squeal_samples[19143]=16447;
squeal_samples[19144]=19059;
squeal_samples[19145]=21563;
squeal_samples[19146]=23944;
squeal_samples[19147]=26236;
squeal_samples[19148]=28419;
squeal_samples[19149]=30500;
squeal_samples[19150]=32501;
squeal_samples[19151]=34401;
squeal_samples[19152]=36224;
squeal_samples[19153]=37962;
squeal_samples[19154]=39625;
squeal_samples[19155]=41208;
squeal_samples[19156]=42723;
squeal_samples[19157]=44172;
squeal_samples[19158]=45550;
squeal_samples[19159]=46877;
squeal_samples[19160]=48132;
squeal_samples[19161]=49344;
squeal_samples[19162]=50485;
squeal_samples[19163]=51593;
squeal_samples[19164]=52643;
squeal_samples[19165]=53173;
squeal_samples[19166]=48825;
squeal_samples[19167]=43497;
squeal_samples[19168]=38507;
squeal_samples[19169]=33839;
squeal_samples[19170]=29466;
squeal_samples[19171]=25376;
squeal_samples[19172]=21557;
squeal_samples[19173]=17969;
squeal_samples[19174]=14620;
squeal_samples[19175]=11485;
squeal_samples[19176]=8551;
squeal_samples[19177]=5991;
squeal_samples[19178]=7474;
squeal_samples[19179]=10476;
squeal_samples[19180]=13349;
squeal_samples[19181]=16100;
squeal_samples[19182]=18726;
squeal_samples[19183]=21246;
squeal_samples[19184]=23645;
squeal_samples[19185]=25941;
squeal_samples[19186]=28140;
squeal_samples[19187]=30235;
squeal_samples[19188]=32241;
squeal_samples[19189]=34160;
squeal_samples[19190]=35985;
squeal_samples[19191]=37735;
squeal_samples[19192]=39406;
squeal_samples[19193]=40999;
squeal_samples[19194]=42529;
squeal_samples[19195]=43978;
squeal_samples[19196]=45372;
squeal_samples[19197]=46698;
squeal_samples[19198]=47967;
squeal_samples[19199]=49176;
squeal_samples[19200]=50334;
squeal_samples[19201]=51443;
squeal_samples[19202]=52500;
squeal_samples[19203]=53296;
squeal_samples[19204]=49506;
squeal_samples[19205]=44127;
squeal_samples[19206]=39101;
squeal_samples[19207]=34389;
squeal_samples[19208]=29988;
squeal_samples[19209]=25857;
squeal_samples[19210]=22006;
squeal_samples[19211]=18390;
squeal_samples[19212]=15018;
squeal_samples[19213]=11850;
squeal_samples[19214]=8901;
squeal_samples[19215]=6171;
squeal_samples[19216]=7083;
squeal_samples[19217]=10099;
squeal_samples[19218]=12984;
squeal_samples[19219]=15752;
squeal_samples[19220]=18391;
squeal_samples[19221]=20928;
squeal_samples[19222]=23336;
squeal_samples[19223]=25649;
squeal_samples[19224]=27856;
squeal_samples[19225]=29967;
squeal_samples[19226]=31986;
squeal_samples[19227]=33913;
squeal_samples[19228]=35751;
squeal_samples[19229]=37511;
squeal_samples[19230]=39188;
squeal_samples[19231]=40792;
squeal_samples[19232]=42331;
squeal_samples[19233]=43786;
squeal_samples[19234]=45193;
squeal_samples[19235]=46522;
squeal_samples[19236]=47803;
squeal_samples[19237]=49016;
squeal_samples[19238]=50181;
squeal_samples[19239]=51294;
squeal_samples[19240]=52356;
squeal_samples[19241]=53375;
squeal_samples[19242]=51011;
squeal_samples[19243]=45531;
squeal_samples[19244]=40422;
squeal_samples[19245]=35617;
squeal_samples[19246]=31140;
squeal_samples[19247]=26936;
squeal_samples[19248]=23014;
squeal_samples[19249]=19335;
squeal_samples[19250]=15893;
squeal_samples[19251]=12679;
squeal_samples[19252]=9666;
squeal_samples[19253]=6848;
squeal_samples[19254]=6389;
squeal_samples[19255]=9391;
squeal_samples[19256]=12310;
squeal_samples[19257]=15108;
squeal_samples[19258]=17776;
squeal_samples[19259]=20335;
squeal_samples[19260]=22770;
squeal_samples[19261]=25112;
squeal_samples[19262]=27337;
squeal_samples[19263]=29472;
squeal_samples[19264]=31512;
squeal_samples[19265]=33456;
squeal_samples[19266]=35316;
squeal_samples[19267]=37098;
squeal_samples[19268]=38793;
squeal_samples[19269]=40419;
squeal_samples[19270]=41962;
squeal_samples[19271]=43450;
squeal_samples[19272]=44852;
squeal_samples[19273]=46214;
squeal_samples[19274]=47490;
squeal_samples[19275]=48733;
squeal_samples[19276]=49898;
squeal_samples[19277]=51030;
squeal_samples[19278]=52095;
squeal_samples[19279]=53132;
squeal_samples[19280]=52222;
squeal_samples[19281]=46878;
squeal_samples[19282]=41664;
squeal_samples[19283]=36794;
squeal_samples[19284]=32231;
squeal_samples[19285]=27958;
squeal_samples[19286]=23968;
squeal_samples[19287]=20229;
squeal_samples[19288]=16736;
squeal_samples[19289]=13456;
squeal_samples[19290]=10396;
squeal_samples[19291]=7529;
squeal_samples[19292]=5971;
squeal_samples[19293]=8639;
squeal_samples[19294]=11591;
squeal_samples[19295]=14411;
squeal_samples[19296]=17114;
squeal_samples[19297]=19701;
squeal_samples[19298]=22169;
squeal_samples[19299]=24528;
squeal_samples[19300]=26781;
squeal_samples[19301]=28943;
squeal_samples[19302]=30996;
squeal_samples[19303]=32975;
squeal_samples[19304]=34851;
squeal_samples[19305]=36653;
squeal_samples[19306]=38369;
squeal_samples[19307]=40010;
squeal_samples[19308]=41571;
squeal_samples[19309]=43072;
squeal_samples[19310]=44500;
squeal_samples[19311]=45868;
squeal_samples[19312]=47167;
squeal_samples[19313]=48418;
squeal_samples[19314]=49607;
squeal_samples[19315]=50743;
squeal_samples[19316]=51823;
squeal_samples[19317]=52869;
squeal_samples[19318]=53012;
squeal_samples[19319]=48228;
squeal_samples[19320]=42918;
squeal_samples[19321]=37977;
squeal_samples[19322]=33327;
squeal_samples[19323]=28998;
squeal_samples[19324]=24925;
squeal_samples[19325]=21130;
squeal_samples[19326]=17575;
squeal_samples[19327]=14244;
squeal_samples[19328]=11134;
squeal_samples[19329]=8217;
squeal_samples[19330]=5899;
squeal_samples[19331]=7871;
squeal_samples[19332]=10851;
squeal_samples[19333]=13710;
squeal_samples[19334]=16438;
squeal_samples[19335]=19054;
squeal_samples[19336]=21550;
squeal_samples[19337]=23932;
squeal_samples[19338]=26221;
squeal_samples[19339]=28397;
squeal_samples[19340]=30487;
squeal_samples[19341]=32474;
squeal_samples[19342]=34382;
squeal_samples[19343]=36197;
squeal_samples[19344]=37937;
squeal_samples[19345]=39595;
squeal_samples[19346]=41180;
squeal_samples[19347]=42694;
squeal_samples[19348]=44138;
squeal_samples[19349]=45517;
squeal_samples[19350]=46837;
squeal_samples[19351]=48094;
squeal_samples[19352]=49302;
squeal_samples[19353]=50447;
squeal_samples[19354]=51548;
squeal_samples[19355]=52597;
squeal_samples[19356]=53394;
squeal_samples[19357]=49591;
squeal_samples[19358]=44205;
squeal_samples[19359]=39171;
squeal_samples[19360]=34450;
squeal_samples[19361]=30034;
squeal_samples[19362]=25910;
squeal_samples[19363]=22045;
squeal_samples[19364]=18433;
squeal_samples[19365]=15040;
squeal_samples[19366]=11882;
squeal_samples[19367]=8914;
squeal_samples[19368]=6189;
squeal_samples[19369]=7095;
squeal_samples[19370]=10102;
squeal_samples[19371]=12992;
squeal_samples[19372]=15755;
squeal_samples[19373]=18399;
squeal_samples[19374]=20925;
squeal_samples[19375]=23341;
squeal_samples[19376]=25640;
squeal_samples[19377]=27852;
squeal_samples[19378]=29956;
squeal_samples[19379]=31974;
squeal_samples[19380]=33905;
squeal_samples[19381]=35732;
squeal_samples[19382]=37498;
squeal_samples[19383]=39168;
squeal_samples[19384]=40780;
squeal_samples[19385]=42306;
squeal_samples[19386]=43767;
squeal_samples[19387]=45170;
squeal_samples[19388]=46501;
squeal_samples[19389]=47777;
squeal_samples[19390]=48988;
squeal_samples[19391]=50155;
squeal_samples[19392]=51266;
squeal_samples[19393]=52331;
squeal_samples[19394]=53342;
squeal_samples[19395]=50982;
squeal_samples[19396]=45508;
squeal_samples[19397]=40386;
squeal_samples[19398]=35588;
squeal_samples[19399]=31105;
squeal_samples[19400]=26900;
squeal_samples[19401]=22974;
squeal_samples[19402]=19301;
squeal_samples[19403]=15852;
squeal_samples[19404]=12643;
squeal_samples[19405]=9623;
squeal_samples[19406]=6809;
squeal_samples[19407]=6352;
squeal_samples[19408]=9354;
squeal_samples[19409]=12272;
squeal_samples[19410]=15065;
squeal_samples[19411]=17734;
squeal_samples[19412]=20290;
squeal_samples[19413]=22729;
squeal_samples[19414]=25067;
squeal_samples[19415]=27295;
squeal_samples[19416]=29428;
squeal_samples[19417]=31471;
squeal_samples[19418]=33411;
squeal_samples[19419]=35274;
squeal_samples[19420]=37053;
squeal_samples[19421]=38753;
squeal_samples[19422]=40367;
squeal_samples[19423]=41924;
squeal_samples[19424]=43395;
squeal_samples[19425]=44815;
squeal_samples[19426]=46160;
squeal_samples[19427]=47453;
squeal_samples[19428]=48678;
squeal_samples[19429]=49861;
squeal_samples[19430]=50981;
squeal_samples[19431]=52059;
squeal_samples[19432]=53082;
squeal_samples[19433]=52184;
squeal_samples[19434]=46825;
squeal_samples[19435]=41625;
squeal_samples[19436]=36744;
squeal_samples[19437]=32183;
squeal_samples[19438]=27914;
squeal_samples[19439]=23920;
squeal_samples[19440]=20181;
squeal_samples[19441]=16687;
squeal_samples[19442]=13408;
squeal_samples[19443]=10348;
squeal_samples[19444]=7481;
squeal_samples[19445]=5920;
squeal_samples[19446]=8595;
squeal_samples[19447]=11537;
squeal_samples[19448]=14374;
squeal_samples[19449]=17061;
squeal_samples[19450]=19656;
squeal_samples[19451]=22119;
squeal_samples[19452]=24478;
squeal_samples[19453]=26737;
squeal_samples[19454]=28888;
squeal_samples[19455]=30955;
squeal_samples[19456]=32921;
squeal_samples[19457]=34806;
squeal_samples[19458]=36602;
squeal_samples[19459]=38322;
squeal_samples[19460]=39961;
squeal_samples[19461]=41529;
squeal_samples[19462]=43021;
squeal_samples[19463]=44456;
squeal_samples[19464]=45815;
squeal_samples[19465]=47122;
squeal_samples[19466]=48368;
squeal_samples[19467]=49558;
squeal_samples[19468]=50695;
squeal_samples[19469]=51783;
squeal_samples[19470]=52815;
squeal_samples[19471]=52972;
squeal_samples[19472]=48169;
squeal_samples[19473]=42880;
squeal_samples[19474]=37920;
squeal_samples[19475]=33286;
squeal_samples[19476]=28945;
squeal_samples[19477]=24878;
squeal_samples[19478]=21082;
squeal_samples[19479]=17526;
squeal_samples[19480]=14196;
squeal_samples[19481]=11085;
squeal_samples[19482]=8170;
squeal_samples[19483]=5850;
squeal_samples[19484]=7822;
squeal_samples[19485]=10804;
squeal_samples[19486]=13659;
squeal_samples[19487]=16393;
squeal_samples[19488]=19004;
squeal_samples[19489]=21502;
squeal_samples[19490]=23884;
squeal_samples[19491]=26171;
squeal_samples[19492]=28351;
squeal_samples[19493]=30437;
squeal_samples[19494]=32426;
squeal_samples[19495]=34334;
squeal_samples[19496]=36148;
squeal_samples[19497]=37889;
squeal_samples[19498]=39546;
squeal_samples[19499]=41131;
squeal_samples[19500]=42648;
squeal_samples[19501]=44088;
squeal_samples[19502]=45469;
squeal_samples[19503]=46787;
squeal_samples[19504]=48047;
squeal_samples[19505]=49254;
squeal_samples[19506]=50399;
squeal_samples[19507]=51499;
squeal_samples[19508]=52548;
squeal_samples[19509]=53347;
squeal_samples[19510]=49542;
squeal_samples[19511]=44158;
squeal_samples[19512]=39120;
squeal_samples[19513]=34404;
squeal_samples[19514]=29990;
squeal_samples[19515]=25862;
squeal_samples[19516]=21997;
squeal_samples[19517]=18384;
squeal_samples[19518]=14993;
squeal_samples[19519]=11832;
squeal_samples[19520]=8867;
squeal_samples[19521]=6139;
squeal_samples[19522]=7047;
squeal_samples[19523]=10055;
squeal_samples[19524]=12944;
squeal_samples[19525]=15704;
squeal_samples[19526]=18354;
squeal_samples[19527]=20873;
squeal_samples[19528]=23295;
squeal_samples[19529]=25591;
squeal_samples[19530]=27804;
squeal_samples[19531]=29906;
squeal_samples[19532]=31930;
squeal_samples[19533]=33850;
squeal_samples[19534]=35691;
squeal_samples[19535]=37443;
squeal_samples[19536]=39125;
squeal_samples[19537]=40727;
squeal_samples[19538]=42261;
squeal_samples[19539]=43716;
squeal_samples[19540]=45124;
squeal_samples[19541]=46451;
squeal_samples[19542]=47728;
squeal_samples[19543]=48941;
squeal_samples[19544]=50103;
squeal_samples[19545]=51223;
squeal_samples[19546]=52276;
squeal_samples[19547]=53297;
squeal_samples[19548]=51703;
squeal_samples[19549]=46232;
squeal_samples[19550]=41059;
squeal_samples[19551]=36219;
squeal_samples[19552]=31692;
squeal_samples[19553]=27448;
squeal_samples[19554]=23482;
squeal_samples[19555]=19769;
squeal_samples[19556]=16297;
squeal_samples[19557]=13042;
squeal_samples[19558]=10005;
squeal_samples[19559]=7159;
squeal_samples[19560]=6099;
squeal_samples[19561]=8983;
squeal_samples[19562]=11910;
squeal_samples[19563]=14725;
squeal_samples[19564]=17403;
squeal_samples[19565]=19975;
squeal_samples[19566]=22426;
squeal_samples[19567]=24769;
squeal_samples[19568]=27006;
squeal_samples[19569]=29155;
squeal_samples[19570]=31201;
squeal_samples[19571]=33160;
squeal_samples[19572]=35028;
squeal_samples[19573]=36816;
squeal_samples[19574]=38519;
squeal_samples[19575]=40151;
squeal_samples[19576]=41712;
squeal_samples[19577]=43189;
squeal_samples[19578]=44616;
squeal_samples[19579]=45969;
squeal_samples[19580]=47268;
squeal_samples[19581]=48501;
squeal_samples[19582]=49685;
squeal_samples[19583]=50815;
squeal_samples[19584]=51894;
squeal_samples[19585]=52925;
squeal_samples[19586]=53069;
squeal_samples[19587]=48267;
squeal_samples[19588]=42964;
squeal_samples[19589]=38002;
squeal_samples[19590]=33349;
squeal_samples[19591]=29009;
squeal_samples[19592]=24932;
squeal_samples[19593]=21135;
squeal_samples[19594]=17568;
squeal_samples[19595]=14240;
squeal_samples[19596]=11115;
squeal_samples[19597]=8202;
squeal_samples[19598]=5871;
squeal_samples[19599]=7841;
squeal_samples[19600]=10827;
squeal_samples[19601]=13678;
squeal_samples[19602]=16404;
squeal_samples[19603]=19017;
squeal_samples[19604]=21514;
squeal_samples[19605]=23892;
squeal_samples[19606]=26176;
squeal_samples[19607]=28356;
squeal_samples[19608]=30434;
squeal_samples[19609]=32433;
squeal_samples[19610]=34326;
squeal_samples[19611]=36147;
squeal_samples[19612]=37884;
squeal_samples[19613]=39536;
squeal_samples[19614]=41125;
squeal_samples[19615]=42635;
squeal_samples[19616]=44080;
squeal_samples[19617]=45461;
squeal_samples[19618]=46775;
squeal_samples[19619]=48041;
squeal_samples[19620]=49237;
squeal_samples[19621]=50384;
squeal_samples[19622]=51484;
squeal_samples[19623]=52533;
squeal_samples[19624]=53484;
squeal_samples[19625]=50337;
squeal_samples[19626]=44898;
squeal_samples[19627]=39813;
squeal_samples[19628]=35048;
squeal_samples[19629]=30595;
squeal_samples[19630]=26416;
squeal_samples[19631]=22526;
squeal_samples[19632]=18865;
squeal_samples[19633]=15453;
squeal_samples[19634]=12250;
squeal_samples[19635]=9262;
squeal_samples[19636]=6461;
squeal_samples[19637]=6683;
squeal_samples[19638]=9712;
squeal_samples[19639]=12608;
squeal_samples[19640]=15387;
squeal_samples[19641]=18035;
squeal_samples[19642]=20581;
squeal_samples[19643]=23005;
squeal_samples[19644]=25318;
squeal_samples[19645]=27539;
squeal_samples[19646]=29654;
squeal_samples[19647]=31679;
squeal_samples[19648]=33617;
squeal_samples[19649]=35461;
squeal_samples[19650]=37231;
squeal_samples[19651]=38918;
squeal_samples[19652]=40525;
squeal_samples[19653]=42064;
squeal_samples[19654]=43539;
squeal_samples[19655]=44934;
squeal_samples[19656]=46279;
squeal_samples[19657]=47560;
squeal_samples[19658]=48779;
squeal_samples[19659]=49949;
squeal_samples[19660]=51069;
squeal_samples[19661]=52134;
squeal_samples[19662]=53156;
squeal_samples[19663]=52244;
squeal_samples[19664]=46883;
squeal_samples[19665]=41671;
squeal_samples[19666]=36786;
squeal_samples[19667]=32219;
squeal_samples[19668]=27941;
squeal_samples[19669]=23937;
squeal_samples[19670]=20196;
squeal_samples[19671]=16696;
squeal_samples[19672]=13411;
squeal_samples[19673]=10347;
squeal_samples[19674]=7478;
squeal_samples[19675]=5908;
squeal_samples[19676]=8580;
squeal_samples[19677]=11523;
squeal_samples[19678]=14351;
squeal_samples[19679]=17047;
squeal_samples[19680]=19629;
squeal_samples[19681]=22097;
squeal_samples[19682]=24450;
squeal_samples[19683]=26705;
squeal_samples[19684]=28863;
squeal_samples[19685]=30922;
squeal_samples[19686]=32890;
squeal_samples[19687]=34769;
squeal_samples[19688]=36568;
squeal_samples[19689]=38283;
squeal_samples[19690]=39920;
squeal_samples[19691]=41485;
squeal_samples[19692]=42981;
squeal_samples[19693]=44408;
squeal_samples[19694]=45773;
squeal_samples[19695]=47075;
squeal_samples[19696]=48316;
squeal_samples[19697]=49511;
squeal_samples[19698]=50639;
squeal_samples[19699]=51729;
squeal_samples[19700]=52765;
squeal_samples[19701]=53280;
squeal_samples[19702]=48923;
squeal_samples[19703]=43569;
squeal_samples[19704]=38566;
squeal_samples[19705]=33888;
squeal_samples[19706]=29494;
squeal_samples[19707]=25400;
squeal_samples[19708]=21557;
squeal_samples[19709]=17969;
squeal_samples[19710]=14609;
squeal_samples[19711]=11461;
squeal_samples[19712]=8519;
squeal_samples[19713]=5942;
squeal_samples[19714]=7427;
squeal_samples[19715]=10425;
squeal_samples[19716]=13290;
squeal_samples[19717]=16036;
squeal_samples[19718]=18661;
squeal_samples[19719]=21174;
squeal_samples[19720]=23568;
squeal_samples[19721]=25859;
squeal_samples[19722]=28051;
squeal_samples[19723]=30146;
squeal_samples[19724]=32150;
squeal_samples[19725]=34063;
squeal_samples[19726]=35889;
squeal_samples[19727]=37634;
squeal_samples[19728]=39302;
squeal_samples[19729]=40897;
squeal_samples[19730]=42414;
squeal_samples[19731]=43868;
squeal_samples[19732]=45252;
squeal_samples[19733]=46581;
squeal_samples[19734]=47844;
squeal_samples[19735]=49055;
squeal_samples[19736]=50214;
squeal_samples[19737]=51315;
squeal_samples[19738]=52369;
squeal_samples[19739]=53379;
squeal_samples[19740]=51010;
squeal_samples[19741]=45523;
squeal_samples[19742]=40397;
squeal_samples[19743]=35590;
squeal_samples[19744]=31097;
squeal_samples[19745]=26890;
squeal_samples[19746]=22958;
squeal_samples[19747]=19278;
squeal_samples[19748]=15827;
squeal_samples[19749]=12603;
squeal_samples[19750]=9586;
squeal_samples[19751]=6765;
squeal_samples[19752]=6304;
squeal_samples[19753]=9304;
squeal_samples[19754]=12218;
squeal_samples[19755]=15010;
squeal_samples[19756]=17676;
squeal_samples[19757]=20234;
squeal_samples[19758]=22670;
squeal_samples[19759]=25002;
squeal_samples[19760]=27228;
squeal_samples[19761]=29367;
squeal_samples[19762]=31397;
squeal_samples[19763]=33342;
squeal_samples[19764]=35202;
squeal_samples[19765]=36979;
squeal_samples[19766]=38675;
squeal_samples[19767]=40293;
squeal_samples[19768]=41841;
squeal_samples[19769]=43319;
squeal_samples[19770]=44735;
squeal_samples[19771]=46077;
squeal_samples[19772]=47365;
squeal_samples[19773]=48599;
squeal_samples[19774]=49771;
squeal_samples[19775]=50897;
squeal_samples[19776]=51969;
squeal_samples[19777]=52991;
squeal_samples[19778]=52660;
squeal_samples[19779]=47524;
squeal_samples[19780]=42261;
squeal_samples[19781]=37346;
squeal_samples[19782]=32734;
squeal_samples[19783]=28427;
squeal_samples[19784]=24386;
squeal_samples[19785]=20615;
squeal_samples[19786]=17083;
squeal_samples[19787]=13774;
squeal_samples[19788]=10682;
squeal_samples[19789]=7794;
squeal_samples[19790]=5800;
squeal_samples[19791]=8162;
squeal_samples[19792]=11131;
squeal_samples[19793]=13964;
squeal_samples[19794]=16684;
squeal_samples[19795]=19275;
squeal_samples[19796]=21758;
squeal_samples[19797]=24126;
squeal_samples[19798]=26392;
squeal_samples[19799]=28562;
squeal_samples[19800]=30630;
squeal_samples[19801]=32615;
squeal_samples[19802]=34501;
squeal_samples[19803]=36309;
squeal_samples[19804]=38034;
squeal_samples[19805]=39685;
squeal_samples[19806]=41257;
squeal_samples[19807]=42762;
squeal_samples[19808]=44194;
squeal_samples[19809]=45566;
squeal_samples[19810]=46883;
squeal_samples[19811]=48128;
squeal_samples[19812]=49327;
squeal_samples[19813]=50464;
squeal_samples[19814]=51561;
squeal_samples[19815]=52603;
squeal_samples[19816]=53392;
squeal_samples[19817]=49577;
squeal_samples[19818]=44184;
squeal_samples[19819]=39141;
squeal_samples[19820]=34412;
squeal_samples[19821]=29995;
squeal_samples[19822]=25856;
squeal_samples[19823]=21988;
squeal_samples[19824]=18369;
squeal_samples[19825]=14978;
squeal_samples[19826]=11806;
squeal_samples[19827]=8842;
squeal_samples[19828]=6107;
squeal_samples[19829]=7011;
squeal_samples[19830]=10018;
squeal_samples[19831]=12907;
squeal_samples[19832]=15664;
squeal_samples[19833]=18303;
squeal_samples[19834]=20831;
squeal_samples[19835]=23235;
squeal_samples[19836]=25545;
squeal_samples[19837]=27746;
squeal_samples[19838]=29859;
squeal_samples[19839]=31865;
squeal_samples[19840]=33793;
squeal_samples[19841]=35626;
squeal_samples[19842]=37385;
squeal_samples[19843]=39058;
squeal_samples[19844]=40665;
squeal_samples[19845]=42192;
squeal_samples[19846]=43652;
squeal_samples[19847]=45055;
squeal_samples[19848]=46376;
squeal_samples[19849]=47660;
squeal_samples[19850]=48871;
squeal_samples[19851]=50035;
squeal_samples[19852]=51147;
squeal_samples[19853]=52203;
squeal_samples[19854]=53222;
squeal_samples[19855]=51629;
squeal_samples[19856]=46150;
squeal_samples[19857]=40982;
squeal_samples[19858]=36137;
squeal_samples[19859]=31608;
squeal_samples[19860]=27363;
squeal_samples[19861]=23394;
squeal_samples[19862]=19687;
squeal_samples[19863]=16210;
squeal_samples[19864]=12957;
squeal_samples[19865]=9916;
squeal_samples[19866]=7070;
squeal_samples[19867]=6013;
squeal_samples[19868]=8892;
squeal_samples[19869]=11825;
squeal_samples[19870]=14630;
squeal_samples[19871]=17316;
squeal_samples[19872]=19881;
squeal_samples[19873]=22338;
squeal_samples[19874]=24675;
squeal_samples[19875]=26925;
squeal_samples[19876]=29061;
squeal_samples[19877]=31112;
squeal_samples[19878]=33069;
squeal_samples[19879]=34937;
squeal_samples[19880]=36726;
squeal_samples[19881]=38427;
squeal_samples[19882]=40056;
squeal_samples[19883]=41615;
squeal_samples[19884]=43099;
squeal_samples[19885]=44524;
squeal_samples[19886]=45878;
squeal_samples[19887]=47173;
squeal_samples[19888]=48410;
squeal_samples[19889]=49593;
squeal_samples[19890]=50719;
squeal_samples[19891]=51802;
squeal_samples[19892]=52829;
squeal_samples[19893]=53342;
squeal_samples[19894]=48969;
squeal_samples[19895]=43618;
squeal_samples[19896]=38605;
squeal_samples[19897]=33917;
squeal_samples[19898]=29524;
squeal_samples[19899]=25419;
squeal_samples[19900]=21575;
squeal_samples[19901]=17978;
squeal_samples[19902]=14614;
squeal_samples[19903]=11460;
squeal_samples[19904]=8518;
squeal_samples[19905]=5939;
squeal_samples[19906]=7420;
squeal_samples[19907]=10411;
squeal_samples[19908]=13281;
squeal_samples[19909]=16017;
squeal_samples[19910]=18647;
squeal_samples[19911]=21150;
squeal_samples[19912]=23546;
squeal_samples[19913]=25838;
squeal_samples[19914]=28027;
squeal_samples[19915]=30126;
squeal_samples[19916]=32120;
squeal_samples[19917]=34033;
squeal_samples[19918]=35859;
squeal_samples[19919]=37604;
squeal_samples[19920]=39266;
squeal_samples[19921]=40859;
squeal_samples[19922]=42378;
squeal_samples[19923]=43831;
squeal_samples[19924]=45217;
squeal_samples[19925]=46541;
squeal_samples[19926]=47805;
squeal_samples[19927]=49018;
squeal_samples[19928]=50168;
squeal_samples[19929]=51272;
squeal_samples[19930]=52329;
squeal_samples[19931]=53336;
squeal_samples[19932]=51737;
squeal_samples[19933]=46251;
squeal_samples[19934]=41075;
squeal_samples[19935]=36223;
squeal_samples[19936]=31686;
squeal_samples[19937]=27437;
squeal_samples[19938]=23463;
squeal_samples[19939]=19742;
squeal_samples[19940]=16264;
squeal_samples[19941]=13007;
squeal_samples[19942]=9963;
squeal_samples[19943]=7112;
squeal_samples[19944]=6047;
squeal_samples[19945]=8930;
squeal_samples[19946]=11858;
squeal_samples[19947]=14662;
squeal_samples[19948]=17339;
squeal_samples[19949]=19907;
squeal_samples[19950]=22363;
squeal_samples[19951]=24693;
squeal_samples[19952]=26940;
squeal_samples[19953]=29079;
squeal_samples[19954]=31128;
squeal_samples[19955]=33081;
squeal_samples[19956]=34946;
squeal_samples[19957]=36734;
squeal_samples[19958]=38437;
squeal_samples[19959]=40063;
squeal_samples[19960]=41625;
squeal_samples[19961]=43100;
squeal_samples[19962]=44529;
squeal_samples[19963]=45875;
squeal_samples[19964]=47176;
squeal_samples[19965]=48407;
squeal_samples[19966]=49592;
squeal_samples[19967]=50716;
squeal_samples[19968]=51794;
squeal_samples[19969]=52827;
squeal_samples[19970]=53340;
squeal_samples[19971]=48965;
squeal_samples[19972]=43613;
squeal_samples[19973]=38594;
squeal_samples[19974]=33907;
squeal_samples[19975]=29514;
squeal_samples[19976]=25407;
squeal_samples[19977]=21565;
squeal_samples[19978]=17968;
squeal_samples[19979]=14598;
squeal_samples[19980]=11450;
squeal_samples[19981]=8503;
squeal_samples[19982]=5925;
squeal_samples[19983]=7402;
squeal_samples[19984]=10394;
squeal_samples[19985]=13266;
squeal_samples[19986]=16002;
squeal_samples[19987]=18623;
squeal_samples[19988]=21136;
squeal_samples[19989]=23525;
squeal_samples[19990]=25819;
squeal_samples[19991]=28011;
squeal_samples[19992]=30105;
squeal_samples[19993]=32103;
squeal_samples[19994]=34013;
squeal_samples[19995]=35841;
squeal_samples[19996]=37585;
squeal_samples[19997]=39249;
squeal_samples[19998]=40839;
squeal_samples[19999]=42360;
squeal_samples[20000]=43813;
squeal_samples[20001]=45197;
squeal_samples[20002]=46524;
squeal_samples[20003]=47785;
squeal_samples[20004]=48995;
squeal_samples[20005]=50148;
squeal_samples[20006]=51251;
squeal_samples[20007]=52301;
squeal_samples[20008]=53316;
squeal_samples[20009]=51709;
squeal_samples[20010]=46235;
squeal_samples[20011]=41050;
squeal_samples[20012]=36201;
squeal_samples[20013]=31660;
squeal_samples[20014]=27412;
squeal_samples[20015]=23441;
squeal_samples[20016]=19722;
squeal_samples[20017]=16248;
squeal_samples[20018]=12980;
squeal_samples[20019]=9941;
squeal_samples[20020]=7086;
squeal_samples[20021]=6029;
squeal_samples[20022]=8907;
squeal_samples[20023]=11833;
squeal_samples[20024]=14638;
squeal_samples[20025]=17322;
squeal_samples[20026]=19881;
squeal_samples[20027]=22340;
squeal_samples[20028]=24675;
squeal_samples[20029]=26914;
squeal_samples[20030]=29057;
squeal_samples[20031]=31103;
squeal_samples[20032]=33057;
squeal_samples[20033]=34923;
squeal_samples[20034]=36708;
squeal_samples[20035]=38415;
squeal_samples[20036]=40038;
squeal_samples[20037]=41600;
squeal_samples[20038]=43079;
squeal_samples[20039]=44501;
squeal_samples[20040]=45855;
squeal_samples[20041]=47149;
squeal_samples[20042]=48385;
squeal_samples[20043]=49567;
squeal_samples[20044]=50693;
squeal_samples[20045]=51769;
squeal_samples[20046]=52804;
squeal_samples[20047]=53315;
squeal_samples[20048]=48943;
squeal_samples[20049]=43587;
squeal_samples[20050]=38572;
squeal_samples[20051]=33880;
squeal_samples[20052]=29494;
squeal_samples[20053]=25380;
squeal_samples[20054]=21544;
squeal_samples[20055]=17940;
squeal_samples[20056]=14578;
squeal_samples[20057]=11422;
squeal_samples[20058]=8483;
squeal_samples[20059]=5899;
squeal_samples[20060]=7383;
squeal_samples[20061]=10372;
squeal_samples[20062]=13239;
squeal_samples[20063]=15980;
squeal_samples[20064]=18600;
squeal_samples[20065]=21110;
squeal_samples[20066]=23503;
squeal_samples[20067]=25793;
squeal_samples[20068]=27988;
squeal_samples[20069]=30081;
squeal_samples[20070]=32080;
squeal_samples[20071]=33987;
squeal_samples[20072]=35820;
squeal_samples[20073]=37558;
squeal_samples[20074]=39226;
squeal_samples[20075]=40816;
squeal_samples[20076]=42333;
squeal_samples[20077]=43793;
squeal_samples[20078]=45171;
squeal_samples[20079]=46500;
squeal_samples[20080]=47761;
squeal_samples[20081]=48972;
squeal_samples[20082]=50122;
squeal_samples[20083]=51228;
squeal_samples[20084]=52279;
squeal_samples[20085]=53288;
squeal_samples[20086]=51690;
squeal_samples[20087]=46208;
squeal_samples[20088]=41026;
squeal_samples[20089]=36179;
squeal_samples[20090]=31633;
squeal_samples[20091]=27392;
squeal_samples[20092]=23414;
squeal_samples[20093]=19701;
squeal_samples[20094]=16220;
squeal_samples[20095]=12960;
squeal_samples[20096]=9913;
squeal_samples[20097]=7067;
squeal_samples[20098]=6001;
squeal_samples[20099]=8884;
squeal_samples[20100]=11809;
squeal_samples[20101]=14615;
squeal_samples[20102]=17296;
squeal_samples[20103]=19860;
squeal_samples[20104]=22312;
squeal_samples[20105]=24654;
squeal_samples[20106]=26889;
squeal_samples[20107]=29033;
squeal_samples[20108]=31080;
squeal_samples[20109]=33031;
squeal_samples[20110]=34902;
squeal_samples[20111]=36682;
squeal_samples[20112]=38391;
squeal_samples[20113]=40016;
squeal_samples[20114]=41574;
squeal_samples[20115]=43056;
squeal_samples[20116]=44478;
squeal_samples[20117]=45828;
squeal_samples[20118]=47130;
squeal_samples[20119]=48355;
squeal_samples[20120]=49549;
squeal_samples[20121]=50664;
squeal_samples[20122]=51748;
squeal_samples[20123]=52780;
squeal_samples[20124]=53288;
squeal_samples[20125]=48923;
squeal_samples[20126]=43560;
squeal_samples[20127]=38551;
squeal_samples[20128]=33853;
squeal_samples[20129]=29472;
squeal_samples[20130]=25354;
squeal_samples[20131]=21522;
squeal_samples[20132]=17917;
squeal_samples[20133]=14550;
squeal_samples[20134]=11404;
squeal_samples[20135]=8452;
squeal_samples[20136]=5881;
squeal_samples[20137]=7355;
squeal_samples[20138]=10350;
squeal_samples[20139]=13215;
squeal_samples[20140]=15956;
squeal_samples[20141]=18575;
squeal_samples[20142]=21087;
squeal_samples[20143]=23478;
squeal_samples[20144]=25770;
squeal_samples[20145]=27964;
squeal_samples[20146]=30057;
squeal_samples[20147]=32056;
squeal_samples[20148]=33964;
squeal_samples[20149]=35793;
squeal_samples[20150]=37537;
squeal_samples[20151]=39200;
squeal_samples[20152]=40794;
squeal_samples[20153]=42309;
squeal_samples[20154]=43767;
squeal_samples[20155]=45148;
squeal_samples[20156]=46476;
squeal_samples[20157]=47738;
squeal_samples[20158]=48945;
squeal_samples[20159]=50103;
squeal_samples[20160]=51199;
squeal_samples[20161]=52258;
squeal_samples[20162]=53263;
squeal_samples[20163]=51666;
squeal_samples[20164]=46183;
squeal_samples[20165]=41005;
squeal_samples[20166]=36151;
squeal_samples[20167]=31612;
squeal_samples[20168]=27367;
squeal_samples[20169]=23390;
squeal_samples[20170]=19678;
squeal_samples[20171]=16194;
squeal_samples[20172]=12938;
squeal_samples[20173]=9889;
squeal_samples[20174]=7041;
squeal_samples[20175]=5981;
squeal_samples[20176]=8857;
squeal_samples[20177]=11786;
squeal_samples[20178]=14592;
squeal_samples[20179]=17268;
squeal_samples[20180]=19841;
squeal_samples[20181]=22285;
squeal_samples[20182]=24633;
squeal_samples[20183]=26862;
squeal_samples[20184]=29010;
squeal_samples[20185]=31055;
squeal_samples[20186]=33010;
squeal_samples[20187]=34874;
squeal_samples[20188]=36662;
squeal_samples[20189]=38363;
squeal_samples[20190]=39994;
squeal_samples[20191]=41551;
squeal_samples[20192]=43029;
squeal_samples[20193]=44458;
squeal_samples[20194]=45801;
squeal_samples[20195]=47106;
squeal_samples[20196]=48333;
squeal_samples[20197]=49522;
squeal_samples[20198]=50642;
squeal_samples[20199]=51725;
squeal_samples[20200]=52752;
squeal_samples[20201]=53270;
squeal_samples[20202]=48892;
squeal_samples[20203]=43542;
squeal_samples[20204]=38522;
squeal_samples[20205]=33833;
squeal_samples[20206]=29445;
squeal_samples[20207]=25333;
squeal_samples[20208]=21495;
squeal_samples[20209]=17894;
squeal_samples[20210]=14527;
squeal_samples[20211]=11378;
squeal_samples[20212]=8431;
squeal_samples[20213]=5853;
squeal_samples[20214]=7336;
squeal_samples[20215]=10320;
squeal_samples[20216]=13197;
squeal_samples[20217]=15927;
squeal_samples[20218]=18554;
squeal_samples[20219]=21062;
squeal_samples[20220]=23454;
squeal_samples[20221]=25746;
squeal_samples[20222]=27940;
squeal_samples[20223]=30031;
squeal_samples[20224]=32035;
squeal_samples[20225]=33937;
squeal_samples[20226]=35771;
squeal_samples[20227]=37511;
squeal_samples[20228]=39178;
squeal_samples[20229]=40767;
squeal_samples[20230]=42288;
squeal_samples[20231]=43741;
squeal_samples[20232]=45124;
squeal_samples[20233]=46452;
squeal_samples[20234]=47714;
squeal_samples[20235]=48920;
squeal_samples[20236]=50081;
squeal_samples[20237]=51172;
squeal_samples[20238]=52235;
squeal_samples[20239]=53238;
squeal_samples[20240]=52314;
squeal_samples[20241]=46945;
squeal_samples[20242]=41709;
squeal_samples[20243]=36816;
squeal_samples[20244]=32225;
squeal_samples[20245]=27942;
squeal_samples[20246]=23924;
squeal_samples[20247]=20175;
squeal_samples[20248]=16660;
squeal_samples[20249]=13374;
squeal_samples[20250]=10294;
squeal_samples[20251]=7420;
squeal_samples[20252]=5841;
squeal_samples[20253]=8507;
squeal_samples[20254]=11453;
squeal_samples[20255]=14266;
squeal_samples[20256]=16962;
squeal_samples[20257]=19539;
squeal_samples[20258]=22005;
squeal_samples[20259]=24355;
squeal_samples[20260]=26607;
squeal_samples[20261]=28759;
squeal_samples[20262]=30811;
squeal_samples[20263]=32781;
squeal_samples[20264]=34655;
squeal_samples[20265]=36446;
squeal_samples[20266]=38164;
squeal_samples[20267]=39791;
squeal_samples[20268]=41361;
squeal_samples[20269]=42848;
squeal_samples[20270]=44278;
squeal_samples[20271]=45641;
squeal_samples[20272]=46936;
squeal_samples[20273]=48181;
squeal_samples[20274]=49372;
squeal_samples[20275]=50497;
squeal_samples[20276]=51587;
squeal_samples[20277]=52618;
squeal_samples[20278]=53559;
squeal_samples[20279]=50391;
squeal_samples[20280]=44946;
squeal_samples[20281]=39833;
squeal_samples[20282]=35066;
squeal_samples[20283]=30584;
squeal_samples[20284]=26409;
squeal_samples[20285]=22490;
squeal_samples[20286]=18826;
squeal_samples[20287]=15399;
squeal_samples[20288]=12190;
squeal_samples[20289]=9188;
squeal_samples[20290]=6387;
squeal_samples[20291]=6594;
squeal_samples[20292]=9622;
squeal_samples[20293]=12515;
squeal_samples[20294]=15288;
squeal_samples[20295]=17936;
squeal_samples[20296]=20473;
squeal_samples[20297]=22894;
squeal_samples[20298]=25204;
squeal_samples[20299]=27418;
squeal_samples[20300]=29530;
squeal_samples[20301]=31557;
squeal_samples[20302]=33482;
squeal_samples[20303]=35329;
squeal_samples[20304]=37089;
squeal_samples[20305]=38776;
squeal_samples[20306]=40383;
squeal_samples[20307]=41921;
squeal_samples[20308]=43388;
squeal_samples[20309]=44784;
squeal_samples[20310]=46130;
squeal_samples[20311]=47400;
squeal_samples[20312]=48627;
squeal_samples[20313]=49787;
squeal_samples[20314]=50901;
squeal_samples[20315]=51968;
squeal_samples[20316]=52986;
squeal_samples[20317]=53116;
squeal_samples[20318]=48295;
squeal_samples[20319]=42974;
squeal_samples[20320]=37999;
squeal_samples[20321]=33341;
squeal_samples[20322]=28972;
squeal_samples[20323]=24898;
squeal_samples[20324]=21075;
squeal_samples[20325]=17508;
squeal_samples[20326]=14158;
squeal_samples[20327]=11031;
squeal_samples[20328]=8109;
squeal_samples[20329]=5765;
squeal_samples[20330]=7735;
squeal_samples[20331]=10710;
squeal_samples[20332]=13560;
squeal_samples[20333]=16278;
squeal_samples[20334]=18887;
squeal_samples[20335]=21377;
squeal_samples[20336]=23756;
squeal_samples[20337]=26036;
squeal_samples[20338]=28211;
squeal_samples[20339]=30291;
squeal_samples[20340]=32277;
squeal_samples[20341]=34175;
squeal_samples[20342]=35990;
squeal_samples[20343]=37719;
squeal_samples[20344]=39374;
squeal_samples[20345]=40955;
squeal_samples[20346]=42467;
squeal_samples[20347]=43906;
squeal_samples[20348]=45285;
squeal_samples[20349]=46599;
squeal_samples[20350]=47857;
squeal_samples[20351]=49060;
squeal_samples[20352]=50203;
squeal_samples[20353]=51298;
squeal_samples[20354]=52342;
squeal_samples[20355]=53347;
squeal_samples[20356]=51738;
squeal_samples[20357]=46251;
squeal_samples[20358]=41060;
squeal_samples[20359]=36203;
squeal_samples[20360]=31652;
squeal_samples[20361]=27408;
squeal_samples[20362]=23412;
squeal_samples[20363]=19703;
squeal_samples[20364]=16207;
squeal_samples[20365]=12955;
squeal_samples[20366]=9899;
squeal_samples[20367]=7046;
squeal_samples[20368]=5980;
squeal_samples[20369]=8851;
squeal_samples[20370]=11781;
squeal_samples[20371]=14583;
squeal_samples[20372]=17262;
squeal_samples[20373]=19823;
squeal_samples[20374]=22274;
squeal_samples[20375]=24612;
squeal_samples[20376]=26848;
squeal_samples[20377]=28987;
squeal_samples[20378]=31032;
squeal_samples[20379]=32987;
squeal_samples[20380]=34853;
squeal_samples[20381]=36634;
squeal_samples[20382]=38336;
squeal_samples[20383]=39966;
squeal_samples[20384]=41516;
squeal_samples[20385]=43004;
squeal_samples[20386]=44421;
squeal_samples[20387]=45771;
squeal_samples[20388]=47067;
squeal_samples[20389]=48299;
squeal_samples[20390]=49484;
squeal_samples[20391]=50603;
squeal_samples[20392]=51684;
squeal_samples[20393]=52712;
squeal_samples[20394]=53486;
squeal_samples[20395]=49659;
squeal_samples[20396]=44246;
squeal_samples[20397]=39189;
squeal_samples[20398]=34449;
squeal_samples[20399]=30015;
squeal_samples[20400]=25865;
squeal_samples[20401]=21988;
squeal_samples[20402]=18351;
squeal_samples[20403]=14948;
squeal_samples[20404]=11775;
squeal_samples[20405]=8793;
squeal_samples[20406]=6057;
squeal_samples[20407]=6946;
squeal_samples[20408]=9953;
squeal_samples[20409]=12834;
squeal_samples[20410]=15587;
squeal_samples[20411]=18223;
squeal_samples[20412]=20743;
squeal_samples[20413]=23154;
squeal_samples[20414]=25449;
squeal_samples[20415]=27653;
squeal_samples[20416]=29755;
squeal_samples[20417]=31766;
squeal_samples[20418]=33682;
squeal_samples[20419]=35524;
squeal_samples[20420]=37267;
squeal_samples[20421]=38948;
squeal_samples[20422]=40541;
squeal_samples[20423]=42072;
squeal_samples[20424]=43527;
squeal_samples[20425]=44926;
squeal_samples[20426]=46252;
squeal_samples[20427]=47527;
squeal_samples[20428]=48733;
squeal_samples[20429]=49900;
squeal_samples[20430]=51006;
squeal_samples[20431]=52063;
squeal_samples[20432]=53076;
squeal_samples[20433]=52731;
squeal_samples[20434]=47579;
squeal_samples[20435]=42304;
squeal_samples[20436]=37360;
squeal_samples[20437]=32740;
squeal_samples[20438]=28414;
squeal_samples[20439]=24368;
squeal_samples[20440]=20578;
squeal_samples[20441]=17042;
squeal_samples[20442]=13720;
squeal_samples[20443]=10622;
squeal_samples[20444]=7716;
squeal_samples[20445]=5717;
squeal_samples[20446]=8076;
squeal_samples[20447]=11040;
squeal_samples[20448]=13870;
squeal_samples[20449]=16581;
squeal_samples[20450]=19169;
squeal_samples[20451]=21645;
squeal_samples[20452]=24015;
squeal_samples[20453]=26274;
squeal_samples[20454]=28444;
squeal_samples[20455]=30508;
squeal_samples[20456]=32484;
squeal_samples[20457]=34370;
squeal_samples[20458]=36174;
squeal_samples[20459]=37896;
squeal_samples[20460]=39538;
squeal_samples[20461]=41115;
squeal_samples[20462]=42607;
squeal_samples[20463]=44054;
squeal_samples[20464]=45414;
squeal_samples[20465]=46727;
squeal_samples[20466]=47973;
squeal_samples[20467]=49164;
squeal_samples[20468]=50303;
squeal_samples[20469]=51399;
squeal_samples[20470]=52436;
squeal_samples[20471]=53430;
squeal_samples[20472]=51046;
squeal_samples[20473]=45545;
squeal_samples[20474]=40402;
squeal_samples[20475]=35581;
squeal_samples[20476]=31074;
squeal_samples[20477]=26847;
squeal_samples[20478]=22914;
squeal_samples[20479]=19212;
squeal_samples[20480]=15761;
squeal_samples[20481]=12516;
squeal_samples[20482]=9497;
squeal_samples[20483]=6666;
squeal_samples[20484]=6194;
squeal_samples[20485]=9191;
squeal_samples[20486]=12102;
squeal_samples[20487]=14886;
squeal_samples[20488]=17549;
squeal_samples[20489]=20100;
squeal_samples[20490]=22533;
squeal_samples[20491]=24859;
squeal_samples[20492]=27090;
squeal_samples[20493]=29215;
squeal_samples[20494]=31248;
squeal_samples[20495]=33188;
squeal_samples[20496]=35046;
squeal_samples[20497]=36813;
squeal_samples[20498]=38507;
squeal_samples[20499]=40125;
squeal_samples[20500]=41670;
squeal_samples[20501]=43149;
squeal_samples[20502]=44555;
squeal_samples[20503]=45902;
squeal_samples[20504]=47181;
squeal_samples[20505]=48419;
squeal_samples[20506]=49581;
squeal_samples[20507]=50708;
squeal_samples[20508]=51776;
squeal_samples[20509]=52801;
squeal_samples[20510]=53305;
squeal_samples[20511]=48926;
squeal_samples[20512]=43559;
squeal_samples[20513]=38544;
squeal_samples[20514]=33843;
squeal_samples[20515]=29446;
squeal_samples[20516]=25331;
squeal_samples[20517]=21483;
squeal_samples[20518]=17881;
squeal_samples[20519]=14506;
squeal_samples[20520]=11350;
squeal_samples[20521]=8402;
squeal_samples[20522]=5816;
squeal_samples[20523]=7292;
squeal_samples[20524]=10287;
squeal_samples[20525]=13150;
squeal_samples[20526]=15888;
squeal_samples[20527]=18511;
squeal_samples[20528]=21014;
squeal_samples[20529]=23402;
squeal_samples[20530]=25692;
squeal_samples[20531]=27888;
squeal_samples[20532]=29972;
squeal_samples[20533]=31976;
squeal_samples[20534]=33880;
squeal_samples[20535]=35706;
squeal_samples[20536]=37449;
squeal_samples[20537]=39112;
squeal_samples[20538]=40705;
squeal_samples[20539]=42216;
squeal_samples[20540]=43674;
squeal_samples[20541]=45054;
squeal_samples[20542]=46383;
squeal_samples[20543]=47638;
squeal_samples[20544]=48847;
squeal_samples[20545]=50003;
squeal_samples[20546]=51100;
squeal_samples[20547]=52157;
squeal_samples[20548]=53164;
squeal_samples[20549]=52810;
squeal_samples[20550]=47651;
squeal_samples[20551]=42364;
squeal_samples[20552]=37423;
squeal_samples[20553]=32794;
squeal_samples[20554]=28462;
squeal_samples[20555]=24410;
squeal_samples[20556]=20620;
squeal_samples[20557]=17070;
squeal_samples[20558]=13750;
squeal_samples[20559]=10642;
squeal_samples[20560]=7738;
squeal_samples[20561]=5732;
squeal_samples[20562]=8092;
squeal_samples[20563]=11044;
squeal_samples[20564]=13880;
squeal_samples[20565]=16584;
squeal_samples[20566]=19181;
squeal_samples[20567]=21649;
squeal_samples[20568]=24018;
squeal_samples[20569]=26275;
squeal_samples[20570]=28441;
squeal_samples[20571]=30502;
squeal_samples[20572]=32485;
squeal_samples[20573]=34361;
squeal_samples[20574]=36168;
squeal_samples[20575]=37885;
squeal_samples[20576]=39530;
squeal_samples[20577]=41104;
squeal_samples[20578]=42602;
squeal_samples[20579]=44034;
squeal_samples[20580]=45403;
squeal_samples[20581]=46710;
squeal_samples[20582]=47959;
squeal_samples[20583]=49150;
squeal_samples[20584]=50287;
squeal_samples[20585]=51380;
squeal_samples[20586]=52414;
squeal_samples[20587]=53410;
squeal_samples[20588]=51797;
squeal_samples[20589]=46297;
squeal_samples[20590]=41102;
squeal_samples[20591]=36239;
squeal_samples[20592]=31683;
squeal_samples[20593]=27426;
squeal_samples[20594]=23434;
squeal_samples[20595]=19709;
squeal_samples[20596]=16214;
squeal_samples[20597]=12951;
squeal_samples[20598]=9894;
squeal_samples[20599]=7029;
squeal_samples[20600]=5970;
squeal_samples[20601]=8837;
squeal_samples[20602]=11764;
squeal_samples[20603]=14560;
squeal_samples[20604]=17237;
squeal_samples[20605]=19801;
squeal_samples[20606]=22247;
squeal_samples[20607]=24586;
squeal_samples[20608]=26817;
squeal_samples[20609]=28961;
squeal_samples[20610]=30996;
squeal_samples[20611]=32952;
squeal_samples[20612]=34813;
squeal_samples[20613]=36599;
squeal_samples[20614]=38298;
squeal_samples[20615]=39918;
squeal_samples[20616]=41480;
squeal_samples[20617]=42954;
squeal_samples[20618]=44379;
squeal_samples[20619]=45724;
squeal_samples[20620]=47020;
squeal_samples[20621]=48252;
squeal_samples[20622]=49429;
squeal_samples[20623]=50555;
squeal_samples[20624]=51631;
squeal_samples[20625]=52661;
squeal_samples[20626]=53587;
squeal_samples[20627]=50423;
squeal_samples[20628]=44956;
squeal_samples[20629]=39850;
squeal_samples[20630]=35060;
squeal_samples[20631]=30584;
squeal_samples[20632]=26389;
squeal_samples[20633]=22475;
squeal_samples[20634]=18805;
squeal_samples[20635]=15365;
squeal_samples[20636]=12158;
squeal_samples[20637]=9151;
squeal_samples[20638]=6342;
squeal_samples[20639]=6547;
squeal_samples[20640]=9572;
squeal_samples[20641]=12461;
squeal_samples[20642]=15235;
squeal_samples[20643]=17874;
squeal_samples[20644]=20410;
squeal_samples[20645]=22827;
squeal_samples[20646]=25141;
squeal_samples[20647]=27352;
squeal_samples[20648]=29464;
squeal_samples[20649]=31488;
squeal_samples[20650]=33410;
squeal_samples[20651]=35259;
squeal_samples[20652]=37013;
squeal_samples[20653]=38700;
squeal_samples[20654]=40301;
squeal_samples[20655]=41842;
squeal_samples[20656]=43303;
squeal_samples[20657]=44705;
squeal_samples[20658]=46042;
squeal_samples[20659]=47319;
squeal_samples[20660]=48540;
squeal_samples[20661]=49705;
squeal_samples[20662]=50814;
squeal_samples[20663]=51882;
squeal_samples[20664]=52897;
squeal_samples[20665]=53400;
squeal_samples[20666]=49003;
squeal_samples[20667]=43642;
squeal_samples[20668]=38603;
squeal_samples[20669]=33904;
squeal_samples[20670]=29490;
squeal_samples[20671]=25377;
squeal_samples[20672]=21521;
squeal_samples[20673]=17914;
squeal_samples[20674]=14534;
squeal_samples[20675]=11372;
squeal_samples[20676]=8419;
squeal_samples[20677]=5831;
squeal_samples[20678]=7306;
squeal_samples[20679]=10290;
squeal_samples[20680]=13159;
squeal_samples[20681]=15892;
squeal_samples[20682]=18512;
squeal_samples[20683]=21014;
squeal_samples[20684]=23403;
squeal_samples[20685]=25688;
squeal_samples[20686]=27875;
squeal_samples[20687]=29965;
squeal_samples[20688]=31963;
squeal_samples[20689]=33870;
squeal_samples[20690]=35692;
squeal_samples[20691]=37431;
squeal_samples[20692]=39097;
squeal_samples[20693]=40685;
squeal_samples[20694]=42198;
squeal_samples[20695]=43654;
squeal_samples[20696]=45034;
squeal_samples[20697]=46353;
squeal_samples[20698]=47621;
squeal_samples[20699]=48822;
squeal_samples[20700]=49978;
squeal_samples[20701]=51075;
squeal_samples[20702]=52123;
squeal_samples[20703]=53133;
squeal_samples[20704]=52777;
squeal_samples[20705]=47619;
squeal_samples[20706]=42334;
squeal_samples[20707]=37389;
squeal_samples[20708]=32762;
squeal_samples[20709]=28431;
squeal_samples[20710]=24371;
squeal_samples[20711]=20586;
squeal_samples[20712]=17029;
squeal_samples[20713]=13713;
squeal_samples[20714]=10607;
squeal_samples[20715]=7696;
squeal_samples[20716]=5695;
squeal_samples[20717]=8048;
squeal_samples[20718]=11013;
squeal_samples[20719]=13837;
squeal_samples[20720]=16545;
squeal_samples[20721]=19134;
squeal_samples[20722]=21611;
squeal_samples[20723]=23970;
squeal_samples[20724]=26238;
squeal_samples[20725]=28391;
squeal_samples[20726]=30467;
squeal_samples[20727]=32435;
squeal_samples[20728]=34324;
squeal_samples[20729]=36121;
squeal_samples[20730]=37844;
squeal_samples[20731]=39487;
squeal_samples[20732]=41056;
squeal_samples[20733]=42559;
squeal_samples[20734]=43991;
squeal_samples[20735]=45361;
squeal_samples[20736]=46659;
squeal_samples[20737]=47915;
squeal_samples[20738]=49102;
squeal_samples[20739]=50245;
squeal_samples[20740]=51326;
squeal_samples[20741]=52370;
squeal_samples[20742]=53365;
squeal_samples[20743]=51755;
squeal_samples[20744]=46253;
squeal_samples[20745]=41056;
squeal_samples[20746]=36189;
squeal_samples[20747]=31636;
squeal_samples[20748]=27376;
squeal_samples[20749]=23388;
squeal_samples[20750]=19665;
squeal_samples[20751]=16172;
squeal_samples[20752]=12902;
squeal_samples[20753]=9849;
squeal_samples[20754]=6991;
squeal_samples[20755]=5918;
squeal_samples[20756]=8792;
squeal_samples[20757]=11712;
squeal_samples[20758]=14514;
squeal_samples[20759]=17187;
squeal_samples[20760]=19755;
squeal_samples[20761]=22199;
squeal_samples[20762]=24536;
squeal_samples[20763]=26769;
squeal_samples[20764]=28913;
squeal_samples[20765]=30947;
squeal_samples[20766]=32907;
squeal_samples[20767]=34762;
squeal_samples[20768]=36552;
squeal_samples[20769]=38248;
squeal_samples[20770]=39879;
squeal_samples[20771]=41426;
squeal_samples[20772]=42914;
squeal_samples[20773]=44323;
squeal_samples[20774]=45682;
squeal_samples[20775]=46967;
squeal_samples[20776]=48206;
squeal_samples[20777]=49380;
squeal_samples[20778]=50508;
squeal_samples[20779]=51582;
squeal_samples[20780]=52613;
squeal_samples[20781]=53539;
squeal_samples[20782]=50374;
squeal_samples[20783]=44909;
squeal_samples[20784]=39800;
squeal_samples[20785]=35014;
squeal_samples[20786]=30535;
squeal_samples[20787]=26341;
squeal_samples[20788]=22427;
squeal_samples[20789]=18755;
squeal_samples[20790]=15319;
squeal_samples[20791]=12108;
squeal_samples[20792]=9104;
squeal_samples[20793]=6293;
squeal_samples[20794]=6498;
squeal_samples[20795]=9526;
squeal_samples[20796]=12411;
squeal_samples[20797]=15186;
squeal_samples[20798]=17828;
squeal_samples[20799]=20365;
squeal_samples[20800]=22780;
squeal_samples[20801]=25094;
squeal_samples[20802]=27300;
squeal_samples[20803]=29420;
squeal_samples[20804]=31437;
squeal_samples[20805]=33363;
squeal_samples[20806]=35210;
squeal_samples[20807]=36967;
squeal_samples[20808]=38648;
squeal_samples[20809]=40258;
squeal_samples[20810]=41788;
squeal_samples[20811]=43259;
squeal_samples[20812]=44656;
squeal_samples[20813]=45992;
squeal_samples[20814]=47274;
squeal_samples[20815]=48488;
squeal_samples[20816]=49660;
squeal_samples[20817]=50764;
squeal_samples[20818]=51835;
squeal_samples[20819]=52848;
squeal_samples[20820]=53351;
squeal_samples[20821]=48957;
squeal_samples[20822]=43591;
squeal_samples[20823]=38559;
squeal_samples[20824]=33850;
squeal_samples[20825]=29448;
squeal_samples[20826]=25324;
squeal_samples[20827]=21476;
squeal_samples[20828]=17864;
squeal_samples[20829]=14485;
squeal_samples[20830]=11326;
squeal_samples[20831]=8369;
squeal_samples[20832]=5786;
squeal_samples[20833]=7253;
squeal_samples[20834]=10246;
squeal_samples[20835]=13107;
squeal_samples[20836]=15847;
squeal_samples[20837]=18463;
squeal_samples[20838]=20966;
squeal_samples[20839]=23353;
squeal_samples[20840]=25641;
squeal_samples[20841]=27828;
squeal_samples[20842]=29915;
squeal_samples[20843]=31916;
squeal_samples[20844]=33821;
squeal_samples[20845]=35643;
squeal_samples[20846]=37384;
squeal_samples[20847]=39049;
squeal_samples[20848]=40635;
squeal_samples[20849]=42153;
squeal_samples[20850]=43603;
squeal_samples[20851]=44986;
squeal_samples[20852]=46307;
squeal_samples[20853]=47570;
squeal_samples[20854]=48777;
squeal_samples[20855]=49928;
squeal_samples[20856]=51026;
squeal_samples[20857]=52076;
squeal_samples[20858]=53086;
squeal_samples[20859]=52726;
squeal_samples[20860]=47574;
squeal_samples[20861]=42282;
squeal_samples[20862]=37343;
squeal_samples[20863]=32715;
squeal_samples[20864]=28380;
squeal_samples[20865]=24326;
squeal_samples[20866]=20533;
squeal_samples[20867]=16985;
squeal_samples[20868]=13663;
squeal_samples[20869]=10559;
squeal_samples[20870]=7649;
squeal_samples[20871]=5643;
squeal_samples[20872]=8004;
squeal_samples[20873]=10962;
squeal_samples[20874]=13790;
squeal_samples[20875]=16497;
squeal_samples[20876]=19085;
squeal_samples[20877]=21563;
squeal_samples[20878]=23923;
squeal_samples[20879]=26187;
squeal_samples[20880]=28347;
squeal_samples[20881]=30414;
squeal_samples[20882]=32391;
squeal_samples[20883]=34273;
squeal_samples[20884]=36073;
squeal_samples[20885]=37797;
squeal_samples[20886]=39437;
squeal_samples[20887]=41009;
squeal_samples[20888]=42509;
squeal_samples[20889]=43944;
squeal_samples[20890]=45310;
squeal_samples[20891]=46615;
squeal_samples[20892]=47862;
squeal_samples[20893]=49057;
squeal_samples[20894]=50194;
squeal_samples[20895]=51278;
squeal_samples[20896]=52322;
squeal_samples[20897]=53315;
squeal_samples[20898]=52380;
squeal_samples[20899]=46990;
squeal_samples[20900]=41737;
squeal_samples[20901]=36833;
squeal_samples[20902]=32227;
squeal_samples[20903]=27931;
squeal_samples[20904]=23899;
squeal_samples[20905]=20137;
squeal_samples[20906]=16613;
squeal_samples[20907]=13315;
squeal_samples[20908]=10231;
squeal_samples[20909]=7343;
squeal_samples[20910]=5762;
squeal_samples[20911]=8417;
squeal_samples[20912]=11354;
squeal_samples[20913]=14172;
squeal_samples[20914]=16857;
squeal_samples[20915]=19433;
squeal_samples[20916]=21893;
squeal_samples[20917]=24235;
squeal_samples[20918]=26485;
squeal_samples[20919]=28632;
squeal_samples[20920]=30686;
squeal_samples[20921]=32648;
squeal_samples[20922]=34523;
squeal_samples[20923]=36310;
squeal_samples[20924]=38023;
squeal_samples[20925]=39654;
squeal_samples[20926]=41212;
squeal_samples[20927]=42705;
squeal_samples[20928]=44126;
squeal_samples[20929]=45484;
squeal_samples[20930]=46780;
squeal_samples[20931]=48026;
squeal_samples[20932]=49205;
squeal_samples[20933]=50341;
squeal_samples[20934]=51418;
squeal_samples[20935]=52456;
squeal_samples[20936]=53440;
squeal_samples[20937]=51820;
squeal_samples[20938]=46310;
squeal_samples[20939]=41112;
squeal_samples[20940]=36235;
squeal_samples[20941]=31675;
squeal_samples[20942]=27406;
squeal_samples[20943]=23415;
squeal_samples[20944]=19686;
squeal_samples[20945]=16188;
squeal_samples[20946]=12912;
squeal_samples[20947]=9853;
squeal_samples[20948]=6991;
squeal_samples[20949]=5917;
squeal_samples[20950]=8785;
squeal_samples[20951]=11708;
squeal_samples[20952]=14504;
squeal_samples[20953]=17181;
squeal_samples[20954]=19737;
squeal_samples[20955]=22187;
squeal_samples[20956]=24515;
squeal_samples[20957]=26756;
squeal_samples[20958]=28887;
squeal_samples[20959]=30926;
squeal_samples[20960]=32883;
squeal_samples[20961]=34741;
squeal_samples[20962]=36524;
squeal_samples[20963]=38220;
squeal_samples[20964]=39845;
squeal_samples[20965]=41392;
squeal_samples[20966]=42881;
squeal_samples[20967]=44285;
squeal_samples[20968]=45641;
squeal_samples[20969]=46932;
squeal_samples[20970]=48163;
squeal_samples[20971]=49344;
squeal_samples[20972]=50466;
squeal_samples[20973]=51546;
squeal_samples[20974]=52565;
squeal_samples[20975]=53557;
squeal_samples[20976]=51147;
squeal_samples[20977]=45634;
squeal_samples[20978]=40472;
squeal_samples[20979]=35637;
squeal_samples[20980]=31120;
squeal_samples[20981]=26883;
squeal_samples[20982]=22932;
squeal_samples[20983]=19222;
squeal_samples[20984]=15752;
squeal_samples[20985]=12509;
squeal_samples[20986]=9473;
squeal_samples[20987]=6634;
squeal_samples[20988]=6157;
squeal_samples[20989]=9147;
squeal_samples[20990]=12054;
squeal_samples[20991]=14837;
squeal_samples[20992]=17495;
squeal_samples[20993]=20040;
squeal_samples[20994]=22469;
squeal_samples[20995]=24795;
squeal_samples[20996]=27012;
squeal_samples[20997]=29136;
squeal_samples[20998]=31165;
squeal_samples[20999]=33103;
squeal_samples[21000]=34958;
squeal_samples[21001]=36728;
squeal_samples[21002]=38414;
squeal_samples[21003]=40034;
squeal_samples[21004]=41571;
squeal_samples[21005]=43046;
squeal_samples[21006]=44448;
squeal_samples[21007]=45797;
squeal_samples[21008]=47076;
squeal_samples[21009]=48306;
squeal_samples[21010]=49469;
squeal_samples[21011]=50594;
squeal_samples[21012]=51660;
squeal_samples[21013]=52684;
squeal_samples[21014]=53605;
squeal_samples[21015]=50429;
squeal_samples[21016]=44953;
squeal_samples[21017]=39844;
squeal_samples[21018]=35043;
squeal_samples[21019]=30560;
squeal_samples[21020]=26361;
squeal_samples[21021]=22441;
squeal_samples[21022]=18765;
squeal_samples[21023]=15322;
squeal_samples[21024]=12106;
squeal_samples[21025]=9096;
squeal_samples[21026]=6281;
squeal_samples[21027]=6484;
squeal_samples[21028]=9510;
squeal_samples[21029]=12389;
squeal_samples[21030]=15168;
squeal_samples[21031]=17798;
squeal_samples[21032]=20341;
squeal_samples[21033]=22753;
squeal_samples[21034]=25066;
squeal_samples[21035]=27271;
squeal_samples[21036]=29385;
squeal_samples[21037]=31403;
squeal_samples[21038]=33329;
squeal_samples[21039]=35169;
squeal_samples[21040]=36926;
squeal_samples[21041]=38611;
squeal_samples[21042]=40215;
squeal_samples[21043]=41745;
squeal_samples[21044]=43212;
squeal_samples[21045]=44611;
squeal_samples[21046]=45946;
squeal_samples[21047]=47225;
squeal_samples[21048]=48434;
squeal_samples[21049]=49612;
squeal_samples[21050]=50710;
squeal_samples[21051]=51786;
squeal_samples[21052]=52790;
squeal_samples[21053]=53556;
squeal_samples[21054]=49710;
squeal_samples[21055]=44288;
squeal_samples[21056]=39211;
squeal_samples[21057]=34455;
squeal_samples[21058]=30011;
squeal_samples[21059]=25844;
squeal_samples[21060]=21955;
squeal_samples[21061]=18310;
squeal_samples[21062]=14895;
squeal_samples[21063]=11709;
squeal_samples[21064]=8721;
squeal_samples[21065]=5972;
squeal_samples[21066]=6864;
squeal_samples[21067]=9861;
squeal_samples[21068]=12736;
squeal_samples[21069]=15487;
squeal_samples[21070]=18117;
squeal_samples[21071]=20635;
squeal_samples[21072]=23031;
squeal_samples[21073]=25335;
squeal_samples[21074]=27526;
squeal_samples[21075]=29628;
squeal_samples[21076]=31634;
squeal_samples[21077]=33551;
squeal_samples[21078]=35385;
squeal_samples[21079]=37132;
squeal_samples[21080]=38804;
squeal_samples[21081]=40397;
squeal_samples[21082]=41926;
squeal_samples[21083]=43376;
squeal_samples[21084]=44770;
squeal_samples[21085]=46095;
squeal_samples[21086]=47370;
squeal_samples[21087]=48577;
squeal_samples[21088]=49737;
squeal_samples[21089]=50839;
squeal_samples[21090]=51893;
squeal_samples[21091]=52909;
squeal_samples[21092]=53399;
squeal_samples[21093]=49005;
squeal_samples[21094]=43624;
squeal_samples[21095]=38588;
squeal_samples[21096]=33876;
squeal_samples[21097]=29459;
squeal_samples[21098]=25333;
squeal_samples[21099]=21472;
squeal_samples[21100]=17861;
squeal_samples[21101]=14478;
squeal_samples[21102]=11311;
squeal_samples[21103]=8348;
squeal_samples[21104]=5764;
squeal_samples[21105]=7225;
squeal_samples[21106]=10219;
squeal_samples[21107]=13070;
squeal_samples[21108]=15811;
squeal_samples[21109]=18428;
squeal_samples[21110]=20929;
squeal_samples[21111]=23313;
squeal_samples[21112]=25601;
squeal_samples[21113]=27783;
squeal_samples[21114]=29874;
squeal_samples[21115]=31863;
squeal_samples[21116]=33775;
squeal_samples[21117]=35594;
squeal_samples[21118]=37331;
squeal_samples[21119]=38995;
squeal_samples[21120]=40577;
squeal_samples[21121]=42102;
squeal_samples[21122]=43541;
squeal_samples[21123]=44927;
squeal_samples[21124]=46246;
squeal_samples[21125]=47509;
squeal_samples[21126]=48713;
squeal_samples[21127]=49865;
squeal_samples[21128]=50965;
squeal_samples[21129]=52009;
squeal_samples[21130]=53025;
squeal_samples[21131]=53130;
squeal_samples[21132]=48298;
squeal_samples[21133]=42960;
squeal_samples[21134]=37968;
squeal_samples[21135]=33294;
squeal_samples[21136]=28914;
squeal_samples[21137]=24822;
squeal_samples[21138]=20998;
squeal_samples[21139]=17411;
squeal_samples[21140]=14056;
squeal_samples[21141]=10920;
squeal_samples[21142]=7983;
squeal_samples[21143]=5641;
squeal_samples[21144]=7598;
squeal_samples[21145]=10567;
squeal_samples[21146]=13413;
squeal_samples[21147]=16130;
squeal_samples[21148]=18729;
squeal_samples[21149]=21224;
squeal_samples[21150]=23592;
squeal_samples[21151]=25873;
squeal_samples[21152]=28035;
squeal_samples[21153]=30118;
squeal_samples[21154]=32095;
squeal_samples[21155]=33997;
squeal_samples[21156]=35802;
squeal_samples[21157]=37534;
squeal_samples[21158]=39186;
squeal_samples[21159]=40758;
squeal_samples[21160]=42272;
squeal_samples[21161]=43703;
squeal_samples[21162]=45083;
squeal_samples[21163]=46392;
squeal_samples[21164]=47649;
squeal_samples[21165]=48847;
squeal_samples[21166]=49989;
squeal_samples[21167]=51088;
squeal_samples[21168]=52130;
squeal_samples[21169]=53130;
squeal_samples[21170]=52767;
squeal_samples[21171]=47601;
squeal_samples[21172]=42305;
squeal_samples[21173]=37357;
squeal_samples[21174]=32718;
squeal_samples[21175]=28379;
squeal_samples[21176]=24320;
squeal_samples[21177]=20525;
squeal_samples[21178]=16968;
squeal_samples[21179]=13638;
squeal_samples[21180]=10528;
squeal_samples[21181]=7617;
squeal_samples[21182]=5613;
squeal_samples[21183]=7966;
squeal_samples[21184]=10920;
squeal_samples[21185]=13742;
squeal_samples[21186]=16450;
squeal_samples[21187]=19037;
squeal_samples[21188]=21516;
squeal_samples[21189]=23869;
squeal_samples[21190]=26135;
squeal_samples[21191]=28293;
squeal_samples[21192]=30356;
squeal_samples[21193]=32326;
squeal_samples[21194]=34215;
squeal_samples[21195]=36011;
squeal_samples[21196]=37731;
squeal_samples[21197]=39374;
squeal_samples[21198]=40943;
squeal_samples[21199]=42442;
squeal_samples[21200]=43874;
squeal_samples[21201]=45236;
squeal_samples[21202]=46544;
squeal_samples[21203]=47788;
squeal_samples[21204]=48982;
squeal_samples[21205]=50118;
squeal_samples[21206]=51205;
squeal_samples[21207]=52244;
squeal_samples[21208]=53236;
squeal_samples[21209]=52871;
squeal_samples[21210]=47694;
squeal_samples[21211]=42399;
squeal_samples[21212]=37439;
squeal_samples[21213]=32796;
squeal_samples[21214]=28451;
squeal_samples[21215]=24386;
squeal_samples[21216]=20581;
squeal_samples[21217]=17022;
squeal_samples[21218]=13693;
squeal_samples[21219]=10571;
squeal_samples[21220]=7664;
squeal_samples[21221]=5645;
squeal_samples[21222]=8007;
squeal_samples[21223]=10954;
squeal_samples[21224]=13781;
squeal_samples[21225]=16479;
squeal_samples[21226]=19069;
squeal_samples[21227]=21542;
squeal_samples[21228]=23895;
squeal_samples[21229]=26155;
squeal_samples[21230]=28313;
squeal_samples[21231]=30377;
squeal_samples[21232]=32346;
squeal_samples[21233]=34231;
squeal_samples[21234]=36029;
squeal_samples[21235]=37749;
squeal_samples[21236]=39386;
squeal_samples[21237]=40956;
squeal_samples[21238]=42449;
squeal_samples[21239]=43885;
squeal_samples[21240]=45245;
squeal_samples[21241]=46554;
squeal_samples[21242]=47796;
squeal_samples[21243]=48989;
squeal_samples[21244]=50126;
squeal_samples[21245]=51210;
squeal_samples[21246]=52248;
squeal_samples[21247]=53240;
squeal_samples[21248]=52874;
squeal_samples[21249]=47701;
squeal_samples[21250]=42396;
squeal_samples[21251]=37438;
squeal_samples[21252]=32796;
squeal_samples[21253]=28449;
squeal_samples[21254]=24384;
squeal_samples[21255]=20582;
squeal_samples[21256]=17018;
squeal_samples[21257]=13694;
squeal_samples[21258]=10569;
squeal_samples[21259]=7657;
squeal_samples[21260]=5645;
squeal_samples[21261]=7998;
squeal_samples[21262]=10950;
squeal_samples[21263]=13771;
squeal_samples[21264]=16482;
squeal_samples[21265]=19060;
squeal_samples[21266]=21536;
squeal_samples[21267]=23888;
squeal_samples[21268]=26148;
squeal_samples[21269]=28309;
squeal_samples[21270]=30368;
squeal_samples[21271]=32342;
squeal_samples[21272]=34220;
squeal_samples[21273]=36023;
squeal_samples[21274]=37736;
squeal_samples[21275]=39380;
squeal_samples[21276]=40945;
squeal_samples[21277]=42446;
squeal_samples[21278]=43869;
squeal_samples[21279]=45242;
squeal_samples[21280]=46539;
squeal_samples[21281]=47792;
squeal_samples[21282]=48981;
squeal_samples[21283]=50114;
squeal_samples[21284]=51203;
squeal_samples[21285]=52243;
squeal_samples[21286]=53231;
squeal_samples[21287]=52870;
squeal_samples[21288]=47688;
squeal_samples[21289]=42382;
squeal_samples[21290]=37430;
squeal_samples[21291]=32780;
squeal_samples[21292]=28439;
squeal_samples[21293]=24372;
squeal_samples[21294]=20569;
squeal_samples[21295]=17008;
squeal_samples[21296]=13680;
squeal_samples[21297]=10559;
squeal_samples[21298]=7643;
squeal_samples[21299]=5635;
squeal_samples[21300]=7985;
squeal_samples[21301]=10937;
squeal_samples[21302]=13763;
squeal_samples[21303]=16464;
squeal_samples[21304]=19055;
squeal_samples[21305]=21517;
squeal_samples[21306]=23882;
squeal_samples[21307]=26132;
squeal_samples[21308]=28298;
squeal_samples[21309]=30357;
squeal_samples[21310]=32328;
squeal_samples[21311]=34211;
squeal_samples[21312]=36008;
squeal_samples[21313]=37725;
squeal_samples[21314]=39369;
squeal_samples[21315]=40932;
squeal_samples[21316]=42434;
squeal_samples[21317]=43858;
squeal_samples[21318]=45228;
squeal_samples[21319]=46529;
squeal_samples[21320]=47781;
squeal_samples[21321]=48965;
squeal_samples[21322]=50106;
squeal_samples[21323]=51189;
squeal_samples[21324]=52231;
squeal_samples[21325]=53221;
squeal_samples[21326]=52856;
squeal_samples[21327]=47675;
squeal_samples[21328]=42375;
squeal_samples[21329]=37411;
squeal_samples[21330]=32774;
squeal_samples[21331]=28424;
squeal_samples[21332]=24361;
squeal_samples[21333]=20557;
squeal_samples[21334]=16996;
squeal_samples[21335]=13667;
squeal_samples[21336]=10548;
squeal_samples[21337]=7637;
squeal_samples[21338]=5622;
squeal_samples[21339]=7975;
squeal_samples[21340]=10922;
squeal_samples[21341]=13753;
squeal_samples[21342]=16451;
squeal_samples[21343]=19043;
squeal_samples[21344]=21508;
squeal_samples[21345]=23865;
squeal_samples[21346]=26124;
squeal_samples[21347]=28285;
squeal_samples[21348]=30343;
squeal_samples[21349]=32320;
squeal_samples[21350]=34195;
squeal_samples[21351]=35998;
squeal_samples[21352]=37714;
squeal_samples[21353]=39354;
squeal_samples[21354]=40923;
squeal_samples[21355]=42420;
squeal_samples[21356]=43847;
squeal_samples[21357]=45216;
squeal_samples[21358]=46516;
squeal_samples[21359]=47769;
squeal_samples[21360]=48955;
squeal_samples[21361]=50092;
squeal_samples[21362]=51179;
squeal_samples[21363]=52217;
squeal_samples[21364]=53210;
squeal_samples[21365]=52844;
squeal_samples[21366]=47664;
squeal_samples[21367]=42360;
squeal_samples[21368]=37405;
squeal_samples[21369]=32754;
squeal_samples[21370]=28420;
squeal_samples[21371]=24343;
squeal_samples[21372]=20548;
squeal_samples[21373]=16983;
squeal_samples[21374]=13656;
squeal_samples[21375]=10534;
squeal_samples[21376]=7628;
squeal_samples[21377]=5606;
squeal_samples[21378]=7966;
squeal_samples[21379]=10909;
squeal_samples[21380]=13741;
squeal_samples[21381]=16441;
squeal_samples[21382]=19028;
squeal_samples[21383]=21496;
squeal_samples[21384]=23856;
squeal_samples[21385]=26109;
squeal_samples[21386]=28274;
squeal_samples[21387]=30333;
squeal_samples[21388]=32304;
squeal_samples[21389]=34187;
squeal_samples[21390]=35984;
squeal_samples[21391]=37702;
squeal_samples[21392]=39343;
squeal_samples[21393]=40911;
squeal_samples[21394]=42407;
squeal_samples[21395]=43837;
squeal_samples[21396]=45202;
squeal_samples[21397]=46507;
squeal_samples[21398]=47754;
squeal_samples[21399]=48945;
squeal_samples[21400]=50079;
squeal_samples[21401]=51166;
squeal_samples[21402]=52208;
squeal_samples[21403]=53195;
squeal_samples[21404]=52835;
squeal_samples[21405]=47649;
squeal_samples[21406]=42351;
squeal_samples[21407]=37390;
squeal_samples[21408]=32745;
squeal_samples[21409]=28406;
squeal_samples[21410]=24331;
squeal_samples[21411]=20539;
squeal_samples[21412]=16967;
squeal_samples[21413]=13647;
squeal_samples[21414]=10522;
squeal_samples[21415]=7613;
squeal_samples[21416]=5600;
squeal_samples[21417]=7947;
squeal_samples[21418]=10904;
squeal_samples[21419]=13723;
squeal_samples[21420]=16433;
squeal_samples[21421]=19013;
squeal_samples[21422]=21488;
squeal_samples[21423]=23840;
squeal_samples[21424]=26101;
squeal_samples[21425]=28259;
squeal_samples[21426]=30321;
squeal_samples[21427]=32294;
squeal_samples[21428]=34174;
squeal_samples[21429]=35972;
squeal_samples[21430]=37690;
squeal_samples[21431]=39332;
squeal_samples[21432]=40897;
squeal_samples[21433]=42398;
squeal_samples[21434]=43822;
squeal_samples[21435]=45191;
squeal_samples[21436]=46495;
squeal_samples[21437]=47743;
squeal_samples[21438]=48932;
squeal_samples[21439]=50068;
squeal_samples[21440]=51154;
squeal_samples[21441]=52194;
squeal_samples[21442]=53187;
squeal_samples[21443]=52818;
squeal_samples[21444]=47642;
squeal_samples[21445]=42336;
squeal_samples[21446]=37379;
squeal_samples[21447]=32735;
squeal_samples[21448]=28389;
squeal_samples[21449]=24325;
squeal_samples[21450]=20521;
squeal_samples[21451]=16962;
squeal_samples[21452]=13628;
squeal_samples[21453]=10516;
squeal_samples[21454]=7597;
squeal_samples[21455]=5589;
squeal_samples[21456]=7937;
squeal_samples[21457]=10888;
squeal_samples[21458]=13716;
squeal_samples[21459]=16418;
squeal_samples[21460]=19003;
squeal_samples[21461]=21475;
squeal_samples[21462]=23827;
squeal_samples[21463]=26092;
squeal_samples[21464]=28243;
squeal_samples[21465]=30315;
squeal_samples[21466]=32276;
squeal_samples[21467]=34167;
squeal_samples[21468]=35956;
squeal_samples[21469]=37682;
squeal_samples[21470]=39316;
squeal_samples[21471]=40889;
squeal_samples[21472]=42382;
squeal_samples[21473]=43814;
squeal_samples[21474]=45177;
squeal_samples[21475]=46485;
squeal_samples[21476]=47728;
squeal_samples[21477]=48923;
squeal_samples[21478]=50054;
squeal_samples[21479]=51143;
squeal_samples[21480]=52184;
squeal_samples[21481]=53171;
squeal_samples[21482]=52810;
squeal_samples[21483]=47627;
squeal_samples[21484]=42326;
squeal_samples[21485]=37367;
squeal_samples[21486]=32722;
squeal_samples[21487]=28378;
squeal_samples[21488]=24313;
squeal_samples[21489]=20508;
squeal_samples[21490]=16951;
squeal_samples[21491]=13617;
squeal_samples[21492]=10502;
squeal_samples[21493]=7587;
squeal_samples[21494]=5576;
squeal_samples[21495]=7925;
squeal_samples[21496]=10878;
squeal_samples[21497]=13701;
squeal_samples[21498]=16408;
squeal_samples[21499]=18991;
squeal_samples[21500]=21461;
squeal_samples[21501]=23820;
squeal_samples[21502]=26073;
squeal_samples[21503]=28239;
squeal_samples[21504]=30297;
squeal_samples[21505]=32266;
squeal_samples[21506]=34156;
squeal_samples[21507]=35942;
squeal_samples[21508]=37674;
squeal_samples[21509]=39300;
squeal_samples[21510]=40879;
squeal_samples[21511]=42370;
squeal_samples[21512]=43801;
squeal_samples[21513]=45168;
squeal_samples[21514]=46469;
squeal_samples[21515]=47720;
squeal_samples[21516]=48907;
squeal_samples[21517]=50046;
squeal_samples[21518]=51129;
squeal_samples[21519]=52172;
squeal_samples[21520]=53160;
squeal_samples[21521]=52797;
squeal_samples[21522]=47616;
squeal_samples[21523]=42314;
squeal_samples[21524]=37353;
squeal_samples[21525]=32713;
squeal_samples[21526]=28364;
squeal_samples[21527]=24302;
squeal_samples[21528]=20497;
squeal_samples[21529]=16937;
squeal_samples[21530]=13606;
squeal_samples[21531]=10489;
squeal_samples[21532]=7577;
squeal_samples[21533]=5562;
squeal_samples[21534]=7916;
squeal_samples[21535]=10863;
squeal_samples[21536]=13690;
squeal_samples[21537]=16396;
squeal_samples[21538]=18979;
squeal_samples[21539]=21451;
squeal_samples[21540]=23805;
squeal_samples[21541]=26063;
squeal_samples[21542]=28226;
squeal_samples[21543]=30284;
squeal_samples[21544]=32258;
squeal_samples[21545]=34139;
squeal_samples[21546]=35934;
squeal_samples[21547]=37657;
squeal_samples[21548]=39294;
squeal_samples[21549]=40862;
squeal_samples[21550]=42361;
squeal_samples[21551]=43788;
squeal_samples[21552]=45154;
squeal_samples[21553]=46459;
squeal_samples[21554]=47707;
squeal_samples[21555]=48896;
squeal_samples[21556]=50033;
squeal_samples[21557]=51116;
squeal_samples[21558]=52160;
squeal_samples[21559]=53147;
squeal_samples[21560]=53254;
squeal_samples[21561]=48395;
squeal_samples[21562]=43052;
squeal_samples[21563]=38043;
squeal_samples[21564]=33355;
squeal_samples[21565]=28970;
squeal_samples[21566]=24856;
squeal_samples[21567]=21024;
squeal_samples[21568]=17425;
squeal_samples[21569]=14060;
squeal_samples[21570]=10919;
squeal_samples[21571]=7970;
squeal_samples[21572]=5623;
squeal_samples[21573]=7574;
squeal_samples[21574]=10539;
squeal_samples[21575]=13378;
squeal_samples[21576]=16097;
squeal_samples[21577]=18689;
squeal_samples[21578]=21179;
squeal_samples[21579]=23541;
squeal_samples[21580]=25816;
squeal_samples[21581]=27983;
squeal_samples[21582]=30057;
squeal_samples[21583]=32034;
squeal_samples[21584]=33924;
squeal_samples[21585]=35736;
squeal_samples[21586]=37458;
squeal_samples[21587]=39108;
squeal_samples[21588]=40684;
squeal_samples[21589]=42189;
squeal_samples[21590]=43627;
squeal_samples[21591]=44994;
squeal_samples[21592]=46312;
squeal_samples[21593]=47558;
squeal_samples[21594]=48760;
squeal_samples[21595]=49901;
squeal_samples[21596]=50991;
squeal_samples[21597]=52033;
squeal_samples[21598]=53026;
squeal_samples[21599]=53512;
squeal_samples[21600]=49097;
squeal_samples[21601]=43702;
squeal_samples[21602]=38650;
squeal_samples[21603]=33919;
squeal_samples[21604]=29501;
squeal_samples[21605]=25354;
squeal_samples[21606]=21486;
squeal_samples[21607]=17862;
squeal_samples[21608]=14468;
squeal_samples[21609]=11291;
squeal_samples[21610]=8324;
squeal_samples[21611]=5724;
squeal_samples[21612]=7187;
squeal_samples[21613]=10175;
squeal_samples[21614]=13023;
squeal_samples[21615]=15758;
squeal_samples[21616]=18365;
squeal_samples[21617]=20858;
squeal_samples[21618]=23248;
squeal_samples[21619]=25528;
squeal_samples[21620]=27712;
squeal_samples[21621]=29796;
squeal_samples[21622]=31788;
squeal_samples[21623]=33685;
squeal_samples[21624]=35506;
squeal_samples[21625]=37240;
squeal_samples[21626]=38903;
squeal_samples[21627]=40478;
squeal_samples[21628]=41998;
squeal_samples[21629]=43440;
squeal_samples[21630]=44825;
squeal_samples[21631]=46140;
squeal_samples[21632]=47401;
squeal_samples[21633]=48600;
squeal_samples[21634]=49748;
squeal_samples[21635]=50844;
squeal_samples[21636]=51894;
squeal_samples[21637]=52898;
squeal_samples[21638]=53643;
squeal_samples[21639]=49788;
squeal_samples[21640]=44346;
squeal_samples[21641]=39254;
squeal_samples[21642]=34481;
squeal_samples[21643]=30027;
squeal_samples[21644]=25848;
squeal_samples[21645]=21944;
squeal_samples[21646]=18294;
squeal_samples[21647]=14864;
squeal_samples[21648]=11675;
squeal_samples[21649]=8666;
squeal_samples[21650]=5923;
squeal_samples[21651]=6792;
squeal_samples[21652]=9793;
squeal_samples[21653]=12665;
squeal_samples[21654]=15409;
squeal_samples[21655]=18038;
squeal_samples[21656]=20543;
squeal_samples[21657]=22946;
squeal_samples[21658]=25237;
squeal_samples[21659]=27426;
squeal_samples[21660]=29533;
squeal_samples[21661]=31526;
squeal_samples[21662]=33446;
squeal_samples[21663]=35267;
squeal_samples[21664]=37019;
squeal_samples[21665]=38684;
squeal_samples[21666]=40277;
squeal_samples[21667]=41800;
squeal_samples[21668]=43251;
squeal_samples[21669]=44643;
squeal_samples[21670]=45967;
squeal_samples[21671]=47230;
squeal_samples[21672]=48443;
squeal_samples[21673]=49599;
squeal_samples[21674]=50702;
squeal_samples[21675]=51758;
squeal_samples[21676]=52764;
squeal_samples[21677]=53677;
squeal_samples[21678]=50480;
squeal_samples[21679]=44994;
squeal_samples[21680]=39858;
squeal_samples[21681]=35054;
squeal_samples[21682]=30555;
squeal_samples[21683]=26343;
squeal_samples[21684]=22410;
squeal_samples[21685]=18725;
squeal_samples[21686]=15269;
squeal_samples[21687]=12044;
squeal_samples[21688]=9023;
squeal_samples[21689]=6200;
squeal_samples[21690]=6405;
squeal_samples[21691]=9412;
squeal_samples[21692]=12304;
squeal_samples[21693]=15057;
squeal_samples[21694]=17701;
squeal_samples[21695]=20230;
squeal_samples[21696]=22639;
squeal_samples[21697]=24947;
squeal_samples[21698]=27151;
squeal_samples[21699]=29256;
squeal_samples[21700]=31276;
squeal_samples[21701]=33195;
squeal_samples[21702]=35037;
squeal_samples[21703]=36788;
squeal_samples[21704]=38470;
squeal_samples[21705]=40073;
squeal_samples[21706]=41600;
squeal_samples[21707]=43064;
squeal_samples[21708]=44455;
squeal_samples[21709]=45793;
squeal_samples[21710]=47066;
squeal_samples[21711]=48285;
squeal_samples[21712]=49445;
squeal_samples[21713]=50555;
squeal_samples[21714]=51616;
squeal_samples[21715]=52626;
squeal_samples[21716]=53600;
squeal_samples[21717]=51179;
squeal_samples[21718]=45651;
squeal_samples[21719]=40471;
squeal_samples[21720]=35628;
squeal_samples[21721]=31089;
squeal_samples[21722]=26838;
squeal_samples[21723]=22873;
squeal_samples[21724]=19156;
squeal_samples[21725]=15677;
squeal_samples[21726]=12424;
squeal_samples[21727]=9380;
squeal_samples[21728]=6531;
squeal_samples[21729]=6049;
squeal_samples[21730]=9032;
squeal_samples[21731]=11938;
squeal_samples[21732]=14710;
squeal_samples[21733]=17368;
squeal_samples[21734]=19907;
squeal_samples[21735]=22336;
squeal_samples[21736]=24647;
squeal_samples[21737]=26868;
squeal_samples[21738]=28989;
squeal_samples[21739]=31014;
squeal_samples[21740]=32951;
squeal_samples[21741]=34796;
squeal_samples[21742]=36565;
squeal_samples[21743]=38253;
squeal_samples[21744]=39864;
squeal_samples[21745]=41401;
squeal_samples[21746]=42870;
squeal_samples[21747]=44276;
squeal_samples[21748]=45618;
squeal_samples[21749]=46897;
squeal_samples[21750]=48121;
squeal_samples[21751]=49288;
squeal_samples[21752]=50405;
squeal_samples[21753]=51475;
squeal_samples[21754]=52488;
squeal_samples[21755]=53467;
squeal_samples[21756]=51834;
squeal_samples[21757]=46305;
squeal_samples[21758]=41084;
squeal_samples[21759]=36205;
squeal_samples[21760]=31625;
squeal_samples[21761]=27348;
squeal_samples[21762]=23342;
squeal_samples[21763]=19596;
squeal_samples[21764]=16089;
squeal_samples[21765]=12806;
squeal_samples[21766]=9740;
squeal_samples[21767]=6861;
squeal_samples[21768]=5787;
squeal_samples[21769]=8647;
squeal_samples[21770]=11563;
squeal_samples[21771]=14361;
squeal_samples[21772]=17027;
squeal_samples[21773]=19582;
squeal_samples[21774]=22026;
squeal_samples[21775]=24351;
squeal_samples[21776]=26586;
squeal_samples[21777]=28717;
squeal_samples[21778]=30751;
squeal_samples[21779]=32702;
squeal_samples[21780]=34561;
squeal_samples[21781]=36337;
squeal_samples[21782]=38034;
squeal_samples[21783]=39653;
squeal_samples[21784]=41201;
squeal_samples[21785]=42683;
squeal_samples[21786]=44089;
squeal_samples[21787]=45443;
squeal_samples[21788]=46730;
squeal_samples[21789]=47959;
squeal_samples[21790]=49137;
squeal_samples[21791]=50257;
squeal_samples[21792]=51333;
squeal_samples[21793]=52350;
squeal_samples[21794]=53337;
squeal_samples[21795]=52380;
squeal_samples[21796]=46972;
squeal_samples[21797]=41712;
squeal_samples[21798]=36778;
squeal_samples[21799]=32175;
squeal_samples[21800]=27853;
squeal_samples[21801]=23814;
squeal_samples[21802]=20042;
squeal_samples[21803]=16503;
squeal_samples[21804]=13194;
squeal_samples[21805]=10096;
squeal_samples[21806]=7203;
squeal_samples[21807]=5613;
squeal_samples[21808]=8263;
squeal_samples[21809]=11196;
squeal_samples[21810]=14004;
squeal_samples[21811]=16690;
squeal_samples[21812]=19262;
squeal_samples[21813]=21713;
squeal_samples[21814]=24055;
squeal_samples[21815]=26300;
squeal_samples[21816]=28445;
squeal_samples[21817]=30491;
squeal_samples[21818]=32450;
squeal_samples[21819]=34322;
squeal_samples[21820]=36106;
squeal_samples[21821]=37813;
squeal_samples[21822]=39443;
squeal_samples[21823]=41003;
squeal_samples[21824]=42489;
squeal_samples[21825]=43904;
squeal_samples[21826]=45265;
squeal_samples[21827]=46556;
squeal_samples[21828]=47800;
squeal_samples[21829]=48981;
squeal_samples[21830]=50105;
squeal_samples[21831]=51191;
squeal_samples[21832]=52212;
squeal_samples[21833]=53205;
squeal_samples[21834]=52830;
squeal_samples[21835]=47647;
squeal_samples[21836]=42337;
squeal_samples[21837]=37368;
squeal_samples[21838]=32719;
squeal_samples[21839]=28368;
squeal_samples[21840]=24294;
squeal_samples[21841]=20482;
squeal_samples[21842]=16924;
squeal_samples[21843]=13583;
squeal_samples[21844]=10462;
squeal_samples[21845]=7543;
squeal_samples[21846]=5526;
squeal_samples[21847]=7880;
squeal_samples[21848]=10824;
squeal_samples[21849]=13648;
squeal_samples[21850]=16351;
squeal_samples[21851]=18931;
squeal_samples[21852]=21400;
squeal_samples[21853]=23754;
squeal_samples[21854]=26011;
squeal_samples[21855]=28169;
squeal_samples[21856]=30227;
squeal_samples[21857]=32201;
squeal_samples[21858]=34076;
squeal_samples[21859]=35879;
squeal_samples[21860]=37592;
squeal_samples[21861]=39233;
squeal_samples[21862]=40793;
squeal_samples[21863]=42295;
squeal_samples[21864]=43717;
squeal_samples[21865]=45090;
squeal_samples[21866]=46388;
squeal_samples[21867]=47635;
squeal_samples[21868]=48821;
squeal_samples[21869]=49960;
squeal_samples[21870]=51043;
squeal_samples[21871]=52081;
squeal_samples[21872]=53068;
squeal_samples[21873]=53542;
squeal_samples[21874]=49122;
squeal_samples[21875]=43723;
squeal_samples[21876]=38664;
squeal_samples[21877]=33929;
squeal_samples[21878]=29498;
squeal_samples[21879]=25354;
squeal_samples[21880]=21478;
squeal_samples[21881]=17844;
squeal_samples[21882]=14450;
squeal_samples[21883]=11274;
squeal_samples[21884]=8294;
squeal_samples[21885]=5696;
squeal_samples[21886]=7159;
squeal_samples[21887]=10138;
squeal_samples[21888]=12986;
squeal_samples[21889]=15718;
squeal_samples[21890]=18322;
squeal_samples[21891]=20825;
squeal_samples[21892]=23196;
squeal_samples[21893]=25487;
squeal_samples[21894]=27661;
squeal_samples[21895]=29744;
squeal_samples[21896]=31739;
squeal_samples[21897]=33634;
squeal_samples[21898]=35456;
squeal_samples[21899]=37184;
squeal_samples[21900]=38846;
squeal_samples[21901]=40425;
squeal_samples[21902]=41938;
squeal_samples[21903]=43383;
squeal_samples[21904]=44759;
squeal_samples[21905]=46082;
squeal_samples[21906]=47332;
squeal_samples[21907]=48541;
squeal_samples[21908]=49684;
squeal_samples[21909]=50784;
squeal_samples[21910]=51826;
squeal_samples[21911]=52830;
squeal_samples[21912]=53734;
squeal_samples[21913]=50536;
squeal_samples[21914]=45042;
squeal_samples[21915]=39895;
squeal_samples[21916]=35085;
squeal_samples[21917]=30577;
squeal_samples[21918]=26363;
squeal_samples[21919]=22423;
squeal_samples[21920]=18727;
squeal_samples[21921]=15276;
squeal_samples[21922]=12042;
squeal_samples[21923]=9018;
squeal_samples[21924]=6188;
squeal_samples[21925]=6388;
squeal_samples[21926]=9396;
squeal_samples[21927]=12281;
squeal_samples[21928]=15035;
squeal_samples[21929]=17679;
squeal_samples[21930]=20201;
squeal_samples[21931]=22612;
squeal_samples[21932]=24914;
squeal_samples[21933]=27118;
squeal_samples[21934]=29223;
squeal_samples[21935]=31236;
squeal_samples[21936]=33164;
squeal_samples[21937]=34995;
squeal_samples[21938]=36754;
squeal_samples[21939]=38423;
squeal_samples[21940]=40030;
squeal_samples[21941]=41556;
squeal_samples[21942]=43019;
squeal_samples[21943]=44412;
squeal_samples[21944]=45748;
squeal_samples[21945]=47017;
squeal_samples[21946]=48235;
squeal_samples[21947]=49391;
squeal_samples[21948]=50505;
squeal_samples[21949]=51559;
squeal_samples[21950]=52578;
squeal_samples[21951]=53543;
squeal_samples[21952]=51903;
squeal_samples[21953]=46373;
squeal_samples[21954]=41137;
squeal_samples[21955]=36248;
squeal_samples[21956]=31666;
squeal_samples[21957]=27380;
squeal_samples[21958]=23363;
squeal_samples[21959]=19620;
squeal_samples[21960]=16104;
squeal_samples[21961]=12818;
squeal_samples[21962]=9746;
squeal_samples[21963]=6867;
squeal_samples[21964]=5782;
squeal_samples[21965]=8647;
squeal_samples[21966]=11560;
squeal_samples[21967]=14352;
squeal_samples[21968]=17019;
squeal_samples[21969]=19572;
squeal_samples[21970]=22009;
squeal_samples[21971]=24337;
squeal_samples[21972]=26568;
squeal_samples[21973]=28696;
squeal_samples[21974]=30731;
squeal_samples[21975]=32679;
squeal_samples[21976]=34537;
squeal_samples[21977]=36306;
squeal_samples[21978]=38006;
squeal_samples[21979]=39622;
squeal_samples[21980]=41174;
squeal_samples[21981]=42646;
squeal_samples[21982]=44059;
squeal_samples[21983]=45405;
squeal_samples[21984]=46691;
squeal_samples[21985]=47924;
squeal_samples[21986]=49097;
squeal_samples[21987]=50215;
squeal_samples[21988]=51293;
squeal_samples[21989]=52315;
squeal_samples[21990]=53296;
squeal_samples[21991]=52914;
squeal_samples[21992]=47719;
squeal_samples[21993]=42402;
squeal_samples[21994]=37432;
squeal_samples[21995]=32772;
squeal_samples[21996]=28415;
squeal_samples[21997]=24338;
squeal_samples[21998]=20520;
squeal_samples[21999]=16956;
squeal_samples[22000]=13607;
squeal_samples[22001]=10485;
squeal_samples[22002]=7556;
squeal_samples[22003]=5543;
squeal_samples[22004]=7882;
squeal_samples[22005]=10833;
squeal_samples[22006]=13651;
squeal_samples[22007]=16348;
squeal_samples[22008]=18933;
squeal_samples[22009]=21396;
squeal_samples[22010]=23753;
squeal_samples[22011]=26007;
squeal_samples[22012]=28164;
squeal_samples[22013]=30218;
squeal_samples[22014]=32187;
squeal_samples[22015]=34065;
squeal_samples[22016]=35866;
squeal_samples[22017]=37577;
squeal_samples[22018]=39212;
squeal_samples[22019]=40780;
squeal_samples[22020]=42273;
squeal_samples[22021]=43697;
squeal_samples[22022]=45065;
squeal_samples[22023]=46363;
squeal_samples[22024]=47608;
squeal_samples[22025]=48799;
squeal_samples[22026]=49929;
squeal_samples[22027]=51018;
squeal_samples[22028]=52049;
squeal_samples[22029]=53042;
squeal_samples[22030]=53509;
squeal_samples[22031]=49092;
squeal_samples[22032]=43692;
squeal_samples[22033]=38627;
squeal_samples[22034]=33898;
squeal_samples[22035]=29467;
squeal_samples[22036]=25318;
squeal_samples[22037]=21441;
squeal_samples[22038]=17809;
squeal_samples[22039]=14412;
squeal_samples[22040]=11233;
squeal_samples[22041]=8257;
squeal_samples[22042]=5661;
squeal_samples[22043]=7116;
squeal_samples[22044]=10098;
squeal_samples[22045]=12948;
squeal_samples[22046]=15677;
squeal_samples[22047]=18281;
squeal_samples[22048]=20781;
squeal_samples[22049]=23163;
squeal_samples[22050]=25443;
squeal_samples[22051]=27619;
squeal_samples[22052]=29704;
squeal_samples[22053]=31689;
squeal_samples[22054]=33595;
squeal_samples[22055]=35407;
squeal_samples[22056]=37142;
squeal_samples[22057]=38801;
squeal_samples[22058]=40380;
squeal_samples[22059]=41894;
squeal_samples[22060]=43338;
squeal_samples[22061]=44721;
squeal_samples[22062]=46031;
squeal_samples[22063]=47294;
squeal_samples[22064]=48490;
squeal_samples[22065]=49640;
squeal_samples[22066]=50735;
squeal_samples[22067]=51786;
squeal_samples[22068]=52787;
squeal_samples[22069]=53693;
squeal_samples[22070]=50489;
squeal_samples[22071]=44993;
squeal_samples[22072]=39850;
squeal_samples[22073]=35037;
squeal_samples[22074]=30536;
squeal_samples[22075]=26316;
squeal_samples[22076]=22374;
squeal_samples[22077]=18681;
squeal_samples[22078]=15229;
squeal_samples[22079]=11995;
squeal_samples[22080]=8970;
squeal_samples[22081]=6142;
squeal_samples[22082]=6340;
squeal_samples[22083]=9350;
squeal_samples[22084]=12237;
squeal_samples[22085]=14991;
squeal_samples[22086]=17628;
squeal_samples[22087]=20157;
squeal_samples[22088]=22570;
squeal_samples[22089]=24865;
squeal_samples[22090]=27073;
squeal_samples[22091]=29180;
squeal_samples[22092]=31189;
squeal_samples[22093]=33119;
squeal_samples[22094]=34946;
squeal_samples[22095]=36706;
squeal_samples[22096]=38379;
squeal_samples[22097]=39979;
squeal_samples[22098]=41514;
squeal_samples[22099]=42967;
squeal_samples[22100]=44367;
squeal_samples[22101]=45701;
squeal_samples[22102]=46969;
squeal_samples[22103]=48190;
squeal_samples[22104]=49346;
squeal_samples[22105]=50460;
squeal_samples[22106]=51512;
squeal_samples[22107]=52530;
squeal_samples[22108]=53497;
squeal_samples[22109]=51855;
squeal_samples[22110]=46326;
squeal_samples[22111]=41091;
squeal_samples[22112]=36200;
squeal_samples[22113]=31620;
squeal_samples[22114]=27331;
squeal_samples[22115]=23323;
squeal_samples[22116]=19573;
squeal_samples[22117]=16055;
squeal_samples[22118]=12775;
squeal_samples[22119]=9693;
squeal_samples[22120]=6825;
squeal_samples[22121]=5732;
squeal_samples[22122]=8601;
squeal_samples[22123]=11513;
squeal_samples[22124]=14305;
squeal_samples[22125]=16972;
squeal_samples[22126]=19524;
squeal_samples[22127]=21961;
squeal_samples[22128]=24292;
squeal_samples[22129]=26520;
squeal_samples[22130]=28649;
squeal_samples[22131]=30684;
squeal_samples[22132]=32632;
squeal_samples[22133]=34488;
squeal_samples[22134]=36262;
squeal_samples[22135]=37956;
squeal_samples[22136]=39578;
squeal_samples[22137]=41124;
squeal_samples[22138]=42602;
squeal_samples[22139]=44008;
squeal_samples[22140]=45363;
squeal_samples[22141]=46639;
squeal_samples[22142]=47882;
squeal_samples[22143]=49044;
squeal_samples[22144]=50174;
squeal_samples[22145]=51242;
squeal_samples[22146]=52270;
squeal_samples[22147]=53248;
squeal_samples[22148]=52867;
squeal_samples[22149]=47671;
squeal_samples[22150]=42358;
squeal_samples[22151]=37380;
squeal_samples[22152]=32730;
squeal_samples[22153]=28364;
squeal_samples[22154]=24292;
squeal_samples[22155]=20475;
squeal_samples[22156]=16905;
squeal_samples[22157]=13563;
squeal_samples[22158]=10437;
squeal_samples[22159]=7508;
squeal_samples[22160]=5497;
squeal_samples[22161]=7835;
squeal_samples[22162]=10785;
squeal_samples[22163]=13605;
squeal_samples[22164]=16301;
squeal_samples[22165]=18885;
squeal_samples[22166]=21350;
squeal_samples[22167]=23706;
squeal_samples[22168]=25958;
squeal_samples[22169]=28120;
squeal_samples[22170]=30169;
squeal_samples[22171]=32140;
squeal_samples[22172]=34020;
squeal_samples[22173]=35816;
squeal_samples[22174]=37532;
squeal_samples[22175]=39164;
squeal_samples[22176]=40732;
squeal_samples[22177]=42227;
squeal_samples[22178]=43652;
squeal_samples[22179]=45015;
squeal_samples[22180]=46317;
squeal_samples[22181]=47562;
squeal_samples[22182]=48747;
squeal_samples[22183]=49890;
squeal_samples[22184]=50964;
squeal_samples[22185]=52006;
squeal_samples[22186]=52994;
squeal_samples[22187]=53460;
squeal_samples[22188]=49048;
squeal_samples[22189]=43642;
squeal_samples[22190]=38582;
squeal_samples[22191]=33850;
squeal_samples[22192]=29421;
squeal_samples[22193]=25268;
squeal_samples[22194]=21398;
squeal_samples[22195]=17757;
squeal_samples[22196]=14371;
squeal_samples[22197]=11180;
squeal_samples[22198]=8214;
squeal_samples[22199]=5611;
squeal_samples[22200]=7072;
squeal_samples[22201]=10047;
squeal_samples[22202]=12905;
squeal_samples[22203]=15625;
squeal_samples[22204]=18239;
squeal_samples[22205]=20731;
squeal_samples[22206]=23117;
squeal_samples[22207]=25395;
squeal_samples[22208]=27572;
squeal_samples[22209]=29657;
squeal_samples[22210]=31642;
squeal_samples[22211]=33549;
squeal_samples[22212]=35357;
squeal_samples[22213]=37099;
squeal_samples[22214]=38748;
squeal_samples[22215]=40339;
squeal_samples[22216]=41842;
squeal_samples[22217]=43295;
squeal_samples[22218]=44670;
squeal_samples[22219]=45987;
squeal_samples[22220]=47243;
squeal_samples[22221]=48447;
squeal_samples[22222]=49588;
squeal_samples[22223]=50692;
squeal_samples[22224]=51735;
squeal_samples[22225]=52741;
squeal_samples[22226]=53694;
squeal_samples[22227]=51266;
squeal_samples[22228]=45720;
squeal_samples[22229]=40522;
squeal_samples[22230]=35672;
squeal_samples[22231]=31115;
squeal_samples[22232]=26863;
squeal_samples[22233]=22874;
squeal_samples[22234]=19156;
squeal_samples[22235]=15664;
squeal_samples[22236]=12400;
squeal_samples[22237]=9345;
squeal_samples[22238]=6494;
squeal_samples[22239]=6001;
squeal_samples[22240]=8985;
squeal_samples[22241]=11879;
squeal_samples[22242]=14650;
squeal_samples[22243]=17306;
squeal_samples[22244]=19841;
squeal_samples[22245]=22263;
squeal_samples[22246]=24576;
squeal_samples[22247]=26789;
squeal_samples[22248]=28907;
squeal_samples[22249]=30930;
squeal_samples[22250]=32862;
squeal_samples[22251]=34709;
squeal_samples[22252]=36470;
squeal_samples[22253]=38154;
squeal_samples[22254]=39764;
squeal_samples[22255]=41302;
squeal_samples[22256]=42764;
squeal_samples[22257]=44174;
squeal_samples[22258]=45504;
squeal_samples[22259]=46790;
squeal_samples[22260]=48007;
squeal_samples[22261]=49180;
squeal_samples[22262]=50288;
squeal_samples[22263]=51358;
squeal_samples[22264]=52373;
squeal_samples[22265]=53344;
squeal_samples[22266]=52962;
squeal_samples[22267]=47754;
squeal_samples[22268]=42435;
squeal_samples[22269]=37451;
squeal_samples[22270]=32788;
squeal_samples[22271]=28426;
squeal_samples[22272]=24338;
squeal_samples[22273]=20524;
squeal_samples[22274]=16945;
squeal_samples[22275]=13598;
squeal_samples[22276]=10467;
squeal_samples[22277]=7532;
squeal_samples[22278]=5515;
squeal_samples[22279]=7855;
squeal_samples[22280]=10804;
squeal_samples[22281]=13623;
squeal_samples[22282]=16315;
squeal_samples[22283]=18897;
squeal_samples[22284]=21360;
squeal_samples[22285]=23711;
squeal_samples[22286]=25965;
squeal_samples[22287]=28117;
squeal_samples[22288]=30176;
squeal_samples[22289]=32140;
squeal_samples[22290]=34017;
squeal_samples[22291]=35815;
squeal_samples[22292]=37521;
squeal_samples[22293]=39164;
squeal_samples[22294]=40721;
squeal_samples[22295]=42221;
squeal_samples[22296]=43640;
squeal_samples[22297]=45010;
squeal_samples[22298]=46301;
squeal_samples[22299]=47548;
squeal_samples[22300]=48736;
squeal_samples[22301]=49866;
squeal_samples[22302]=50953;
squeal_samples[22303]=51985;
squeal_samples[22304]=52980;
squeal_samples[22305]=53707;
squeal_samples[22306]=49839;
squeal_samples[22307]=44376;
squeal_samples[22308]=39275;
squeal_samples[22309]=34488;
squeal_samples[22310]=30015;
squeal_samples[22311]=25826;
squeal_samples[22312]=21914;
squeal_samples[22313]=18246;
squeal_samples[22314]=14814;
squeal_samples[22315]=11606;
squeal_samples[22316]=8599;
squeal_samples[22317]=5837;
squeal_samples[22318]=6710;
squeal_samples[22319]=9704;
squeal_samples[22320]=12567;
squeal_samples[22321]=15312;
squeal_samples[22322]=17926;
squeal_samples[22323]=20439;
squeal_samples[22324]=22830;
squeal_samples[22325]=25122;
squeal_samples[22326]=27308;
squeal_samples[22327]=29404;
squeal_samples[22328]=31402;
squeal_samples[22329]=33310;
squeal_samples[22330]=35135;
squeal_samples[22331]=36882;
squeal_samples[22332]=38541;
squeal_samples[22333]=40138;
squeal_samples[22334]=41652;
squeal_samples[22335]=43105;
squeal_samples[22336]=44491;
squeal_samples[22337]=45814;
squeal_samples[22338]=47079;
squeal_samples[22339]=48284;
squeal_samples[22340]=49437;
squeal_samples[22341]=50537;
squeal_samples[22342]=51596;
squeal_samples[22343]=52599;
squeal_samples[22344]=53561;
squeal_samples[22345]=51913;
squeal_samples[22346]=46369;
squeal_samples[22347]=41139;
squeal_samples[22348]=36234;
squeal_samples[22349]=31648;
squeal_samples[22350]=27354;
squeal_samples[22351]=23332;
squeal_samples[22352]=19584;
squeal_samples[22353]=16061;
squeal_samples[22354]=12772;
squeal_samples[22355]=9692;
squeal_samples[22356]=6809;
squeal_samples[22357]=5725;
squeal_samples[22358]=8581;
squeal_samples[22359]=11500;
squeal_samples[22360]=14280;
squeal_samples[22361]=16952;
squeal_samples[22362]=19496;
squeal_samples[22363]=21933;
squeal_samples[22364]=24266;
squeal_samples[22365]=26485;
squeal_samples[22366]=28619;
squeal_samples[22367]=30649;
squeal_samples[22368]=32595;
squeal_samples[22369]=34448;
squeal_samples[22370]=36226;
squeal_samples[22371]=37916;
squeal_samples[22372]=39535;
squeal_samples[22373]=41081;
squeal_samples[22374]=42556;
squeal_samples[22375]=43969;
squeal_samples[22376]=45313;
squeal_samples[22377]=46601;
squeal_samples[22378]=47828;
squeal_samples[22379]=49000;
squeal_samples[22380]=50119;
squeal_samples[22381]=51192;
squeal_samples[22382]=52212;
squeal_samples[22383]=53195;
squeal_samples[22384]=53284;
squeal_samples[22385]=48416;
squeal_samples[22386]=43045;
squeal_samples[22387]=38026;
squeal_samples[22388]=33315;
squeal_samples[22389]=28924;
squeal_samples[22390]=24797;
squeal_samples[22391]=20951;
squeal_samples[22392]=17343;
squeal_samples[22393]=13970;
squeal_samples[22394]=10811;
squeal_samples[22395]=7858;
squeal_samples[22396]=5500;
squeal_samples[22397]=7444;
squeal_samples[22398]=10412;
squeal_samples[22399]=13236;
squeal_samples[22400]=15953;
squeal_samples[22401]=18545;
squeal_samples[22402]=21019;
squeal_samples[22403]=23392;
squeal_samples[22404]=25648;
squeal_samples[22405]=27821;
squeal_samples[22406]=29887;
squeal_samples[22407]=31869;
squeal_samples[22408]=33752;
squeal_samples[22409]=35556;
squeal_samples[22410]=37284;
squeal_samples[22411]=38922;
squeal_samples[22412]=40503;
squeal_samples[22413]=41994;
squeal_samples[22414]=43437;
squeal_samples[22415]=44802;
squeal_samples[22416]=46112;
squeal_samples[22417]=47358;
squeal_samples[22418]=48556;
squeal_samples[22419]=49693;
squeal_samples[22420]=50784;
squeal_samples[22421]=51823;
squeal_samples[22422]=52825;
squeal_samples[22423]=53715;
squeal_samples[22424]=50510;
squeal_samples[22425]=45004;
squeal_samples[22426]=39860;
squeal_samples[22427]=35031;
squeal_samples[22428]=30525;
squeal_samples[22429]=26300;
squeal_samples[22430]=22357;
squeal_samples[22431]=18656;
squeal_samples[22432]=15197;
squeal_samples[22433]=11962;
squeal_samples[22434]=8926;
squeal_samples[22435]=6100;
squeal_samples[22436]=6288;
squeal_samples[22437]=9303;
squeal_samples[22438]=12177;
squeal_samples[22439]=14940;
squeal_samples[22440]=17573;
squeal_samples[22441]=20097;
squeal_samples[22442]=22508;
squeal_samples[22443]=24804;
squeal_samples[22444]=27007;
squeal_samples[22445]=29115;
squeal_samples[22446]=31120;
squeal_samples[22447]=33044;
squeal_samples[22448]=34876;
squeal_samples[22449]=36629;
squeal_samples[22450]=38308;
squeal_samples[22451]=39903;
squeal_samples[22452]=41436;
squeal_samples[22453]=42888;
squeal_samples[22454]=44289;
squeal_samples[22455]=45616;
squeal_samples[22456]=46884;
squeal_samples[22457]=48105;
squeal_samples[22458]=49258;
squeal_samples[22459]=50368;
squeal_samples[22460]=51429;
squeal_samples[22461]=52439;
squeal_samples[22462]=53405;
squeal_samples[22463]=52442;
squeal_samples[22464]=47015;
squeal_samples[22465]=41737;
squeal_samples[22466]=36794;
squeal_samples[22467]=32169;
squeal_samples[22468]=27841;
squeal_samples[22469]=23785;
squeal_samples[22470]=20005;
squeal_samples[22471]=16455;
squeal_samples[22472]=13139;
squeal_samples[22473]=10030;
squeal_samples[22474]=7131;
squeal_samples[22475]=5521;
squeal_samples[22476]=8176;
squeal_samples[22477]=11101;
squeal_samples[22478]=13907;
squeal_samples[22479]=16589;
squeal_samples[22480]=19151;
squeal_samples[22481]=21600;
squeal_samples[22482]=23942;
squeal_samples[22483]=26181;
squeal_samples[22484]=28320;
squeal_samples[22485]=30366;
squeal_samples[22486]=32319;
squeal_samples[22487]=34189;
squeal_samples[22488]=35969;
squeal_samples[22489]=37679;
squeal_samples[22490]=39299;
squeal_samples[22491]=40860;
squeal_samples[22492]=42341;
squeal_samples[22493]=43759;
squeal_samples[22494]=45110;
squeal_samples[22495]=46408;
squeal_samples[22496]=47640;
squeal_samples[22497]=48820;
squeal_samples[22498]=49947;
squeal_samples[22499]=51025;
squeal_samples[22500]=52054;
squeal_samples[22501]=53036;
squeal_samples[22502]=53508;
squeal_samples[22503]=49073;
squeal_samples[22504]=43664;
squeal_samples[22505]=38597;
squeal_samples[22506]=33851;
squeal_samples[22507]=29421;
squeal_samples[22508]=25261;
squeal_samples[22509]=21382;
squeal_samples[22510]=17749;
squeal_samples[22511]=14341;
squeal_samples[22512]=11162;
squeal_samples[22513]=8181;
squeal_samples[22514]=5574;
squeal_samples[22515]=7028;
squeal_samples[22516]=10012;
squeal_samples[22517]=12853;
squeal_samples[22518]=15587;
squeal_samples[22519]=18187;
squeal_samples[22520]=20684;
squeal_samples[22521]=23063;
squeal_samples[22522]=25341;
squeal_samples[22523]=27516;
squeal_samples[22524]=29599;
squeal_samples[22525]=31588;
squeal_samples[22526]=33483;
squeal_samples[22527]=35300;
squeal_samples[22528]=37035;
squeal_samples[22529]=38688;
squeal_samples[22530]=40270;
squeal_samples[22531]=41781;
squeal_samples[22532]=43222;
squeal_samples[22533]=44598;
squeal_samples[22534]=45919;
squeal_samples[22535]=47171;
squeal_samples[22536]=48373;
squeal_samples[22537]=49517;
squeal_samples[22538]=50617;
squeal_samples[22539]=51658;
squeal_samples[22540]=52662;
squeal_samples[22541]=53620;
squeal_samples[22542]=51968;
squeal_samples[22543]=46415;
squeal_samples[22544]=41175;
squeal_samples[22545]=36264;
squeal_samples[22546]=31675;
squeal_samples[22547]=27376;
squeal_samples[22548]=23350;
squeal_samples[22549]=19594;
squeal_samples[22550]=16068;
squeal_samples[22551]=12774;
squeal_samples[22552]=9690;
squeal_samples[22553]=6807;
squeal_samples[22554]=5713;
squeal_samples[22555]=8572;
squeal_samples[22556]=11483;
squeal_samples[22557]=14266;
squeal_samples[22558]=16936;
squeal_samples[22559]=19480;
squeal_samples[22560]=21919;
squeal_samples[22561]=24243;
squeal_samples[22562]=26465;
squeal_samples[22563]=28593;
squeal_samples[22564]=30622;
squeal_samples[22565]=32568;
squeal_samples[22566]=34424;
squeal_samples[22567]=36192;
squeal_samples[22568]=37885;
squeal_samples[22569]=39504;
squeal_samples[22570]=41047;
squeal_samples[22571]=42520;
squeal_samples[22572]=43931;
squeal_samples[22573]=45276;
squeal_samples[22574]=46559;
squeal_samples[22575]=47788;
squeal_samples[22576]=48960;
squeal_samples[22577]=50074;
squeal_samples[22578]=51150;
squeal_samples[22579]=52169;
squeal_samples[22580]=53149;
squeal_samples[22581]=53609;
squeal_samples[22582]=49169;
squeal_samples[22583]=43754;
squeal_samples[22584]=38681;
squeal_samples[22585]=33931;
squeal_samples[22586]=29490;
squeal_samples[22587]=25324;
squeal_samples[22588]=21440;
squeal_samples[22589]=17799;
squeal_samples[22590]=14390;
squeal_samples[22591]=11203;
squeal_samples[22592]=8217;
squeal_samples[22593]=5609;
squeal_samples[22594]=7066;
squeal_samples[22595]=10039;
squeal_samples[22596]=12889;
squeal_samples[22597]=15607;
squeal_samples[22598]=18215;
squeal_samples[22599]=20709;
squeal_samples[22600]=23077;
squeal_samples[22601]=25361;
squeal_samples[22602]=27534;
squeal_samples[22603]=29616;
squeal_samples[22604]=31599;
squeal_samples[22605]=33496;
squeal_samples[22606]=35306;
squeal_samples[22607]=37038;
squeal_samples[22608]=38693;
squeal_samples[22609]=40272;
squeal_samples[22610]=41785;
squeal_samples[22611]=43227;
squeal_samples[22612]=44599;
squeal_samples[22613]=45919;
squeal_samples[22614]=47168;
squeal_samples[22615]=48372;
squeal_samples[22616]=49516;
squeal_samples[22617]=50608;
squeal_samples[22618]=51656;
squeal_samples[22619]=52657;
squeal_samples[22620]=53610;
squeal_samples[22621]=51957;
squeal_samples[22622]=46407;
squeal_samples[22623]=41161;
squeal_samples[22624]=36259;
squeal_samples[22625]=31661;
squeal_samples[22626]=27363;
squeal_samples[22627]=23339;
squeal_samples[22628]=19578;
squeal_samples[22629]=16060;
squeal_samples[22630]=12755;
squeal_samples[22631]=9678;
squeal_samples[22632]=6785;
squeal_samples[22633]=5701;
squeal_samples[22634]=8556;
squeal_samples[22635]=11466;
squeal_samples[22636]=14252;
squeal_samples[22637]=16915;
squeal_samples[22638]=19463;
squeal_samples[22639]=21901;
squeal_samples[22640]=24223;
squeal_samples[22641]=26450;
squeal_samples[22642]=28572;
squeal_samples[22643]=30605;
squeal_samples[22644]=32551;
squeal_samples[22645]=34398;
squeal_samples[22646]=36175;
squeal_samples[22647]=37867;
squeal_samples[22648]=39485;
squeal_samples[22649]=41024;
squeal_samples[22650]=42504;
squeal_samples[22651]=43903;
squeal_samples[22652]=45257;
squeal_samples[22653]=46536;
squeal_samples[22654]=47770;
squeal_samples[22655]=48936;
squeal_samples[22656]=50061;
squeal_samples[22657]=51128;
squeal_samples[22658]=52153;
squeal_samples[22659]=53126;
squeal_samples[22660]=53588;
squeal_samples[22661]=49153;
squeal_samples[22662]=43730;
squeal_samples[22663]=38657;
squeal_samples[22664]=33910;
squeal_samples[22665]=29467;
squeal_samples[22666]=25311;
squeal_samples[22667]=21417;
squeal_samples[22668]=17780;
squeal_samples[22669]=14364;
squeal_samples[22670]=11180;
squeal_samples[22671]=8194;
squeal_samples[22672]=5584;
squeal_samples[22673]=7044;
squeal_samples[22674]=10015;
squeal_samples[22675]=12865;
squeal_samples[22676]=15584;
squeal_samples[22677]=18193;
squeal_samples[22678]=20682;
squeal_samples[22679]=23062;
squeal_samples[22680]=25336;
squeal_samples[22681]=27511;
squeal_samples[22682]=29593;
squeal_samples[22683]=31575;
squeal_samples[22684]=33472;
squeal_samples[22685]=35283;
squeal_samples[22686]=37020;
squeal_samples[22687]=38669;
squeal_samples[22688]=40254;
squeal_samples[22689]=41763;
squeal_samples[22690]=43199;
squeal_samples[22691]=44582;
squeal_samples[22692]=45889;
squeal_samples[22693]=47150;
squeal_samples[22694]=48344;
squeal_samples[22695]=49494;
squeal_samples[22696]=50590;
squeal_samples[22697]=51634;
squeal_samples[22698]=52630;
squeal_samples[22699]=53590;
squeal_samples[22700]=51935;
squeal_samples[22701]=46387;
squeal_samples[22702]=41137;
squeal_samples[22703]=36234;
squeal_samples[22704]=31639;
squeal_samples[22705]=27337;
squeal_samples[22706]=23317;
squeal_samples[22707]=19556;
squeal_samples[22708]=16033;
squeal_samples[22709]=12736;
squeal_samples[22710]=9650;
squeal_samples[22711]=6770;
squeal_samples[22712]=5676;
squeal_samples[22713]=8533;
squeal_samples[22714]=11443;
squeal_samples[22715]=14228;
squeal_samples[22716]=16891;
squeal_samples[22717]=19440;
squeal_samples[22718]=21878;
squeal_samples[22719]=24199;
squeal_samples[22720]=26427;
squeal_samples[22721]=28547;
squeal_samples[22722]=30583;
squeal_samples[22723]=32526;
squeal_samples[22724]=34376;
squeal_samples[22725]=36151;
squeal_samples[22726]=37843;
squeal_samples[22727]=39462;
squeal_samples[22728]=41001;
squeal_samples[22729]=42477;
squeal_samples[22730]=43886;
squeal_samples[22731]=45225;
squeal_samples[22732]=46522;
squeal_samples[22733]=47737;
squeal_samples[22734]=48922;
squeal_samples[22735]=50029;
squeal_samples[22736]=51110;
squeal_samples[22737]=52125;
squeal_samples[22738]=53107;
squeal_samples[22739]=53562;
squeal_samples[22740]=49130;
squeal_samples[22741]=43706;
squeal_samples[22742]=38633;
squeal_samples[22743]=33888;
squeal_samples[22744]=29443;
squeal_samples[22745]=25285;
squeal_samples[22746]=21397;
squeal_samples[22747]=17754;
squeal_samples[22748]=14342;
squeal_samples[22749]=11156;
squeal_samples[22750]=8169;
squeal_samples[22751]=5563;
squeal_samples[22752]=7018;
squeal_samples[22753]=9994;
squeal_samples[22754]=12839;
squeal_samples[22755]=15563;
squeal_samples[22756]=18165;
squeal_samples[22757]=20663;
squeal_samples[22758]=23036;
squeal_samples[22759]=25314;
squeal_samples[22760]=27487;
squeal_samples[22761]=29567;
squeal_samples[22762]=31555;
squeal_samples[22763]=33446;
squeal_samples[22764]=35262;
squeal_samples[22765]=36994;
squeal_samples[22766]=38646;
squeal_samples[22767]=40232;
squeal_samples[22768]=41737;
squeal_samples[22769]=43180;
squeal_samples[22770]=44552;
squeal_samples[22771]=45872;
squeal_samples[22772]=47121;
squeal_samples[22773]=48324;
squeal_samples[22774]=49469;
squeal_samples[22775]=50567;
squeal_samples[22776]=51610;
squeal_samples[22777]=52607;
squeal_samples[22778]=53566;
squeal_samples[22779]=51912;
squeal_samples[22780]=46363;
squeal_samples[22781]=41113;
squeal_samples[22782]=36212;
squeal_samples[22783]=31613;
squeal_samples[22784]=27318;
squeal_samples[22785]=23288;
squeal_samples[22786]=19536;
squeal_samples[22787]=16007;
squeal_samples[22788]=12716;
squeal_samples[22789]=9623;
squeal_samples[22790]=6749;
squeal_samples[22791]=5650;
squeal_samples[22792]=8510;
squeal_samples[22793]=11421;
squeal_samples[22794]=14202;
squeal_samples[22795]=16870;
squeal_samples[22796]=19416;
squeal_samples[22797]=21852;
squeal_samples[22798]=24179;
squeal_samples[22799]=26400;
squeal_samples[22800]=28526;
squeal_samples[22801]=30559;
squeal_samples[22802]=32502;
squeal_samples[22803]=34353;
squeal_samples[22804]=36128;
squeal_samples[22805]=37818;
squeal_samples[22806]=39439;
squeal_samples[22807]=40977;
squeal_samples[22808]=42455;
squeal_samples[22809]=43860;
squeal_samples[22810]=45207;
squeal_samples[22811]=46490;
squeal_samples[22812]=47722;
squeal_samples[22813]=48889;
squeal_samples[22814]=50015;
squeal_samples[22815]=51080;
squeal_samples[22816]=52107;
squeal_samples[22817]=53078;
squeal_samples[22818]=53541;
squeal_samples[22819]=49106;
squeal_samples[22820]=43683;
squeal_samples[22821]=38610;
squeal_samples[22822]=33862;
squeal_samples[22823]=29423;
squeal_samples[22824]=25258;
squeal_samples[22825]=21378;
squeal_samples[22826]=17724;
squeal_samples[22827]=14325;
squeal_samples[22828]=11126;
squeal_samples[22829]=8152;
squeal_samples[22830]=5534;
squeal_samples[22831]=6998;
squeal_samples[22832]=9969;
squeal_samples[22833]=12816;
squeal_samples[22834]=15538;
squeal_samples[22835]=18145;
squeal_samples[22836]=20635;
squeal_samples[22837]=23017;
squeal_samples[22838]=25287;
squeal_samples[22839]=27465;
squeal_samples[22840]=29545;
squeal_samples[22841]=31528;
squeal_samples[22842]=33425;
squeal_samples[22843]=35236;
squeal_samples[22844]=36974;
squeal_samples[22845]=38620;
squeal_samples[22846]=40210;
squeal_samples[22847]=41712;
squeal_samples[22848]=43156;
squeal_samples[22849]=44531;
squeal_samples[22850]=45846;
squeal_samples[22851]=47100;
squeal_samples[22852]=48298;
squeal_samples[22853]=49447;
squeal_samples[22854]=50542;
squeal_samples[22855]=51589;
squeal_samples[22856]=52581;
squeal_samples[22857]=53545;
squeal_samples[22858]=51885;
squeal_samples[22859]=46342;
squeal_samples[22860]=41088;
squeal_samples[22861]=36190;
squeal_samples[22862]=31589;
squeal_samples[22863]=27294;
squeal_samples[22864]=23265;
squeal_samples[22865]=19512;
squeal_samples[22866]=15984;
squeal_samples[22867]=12691;
squeal_samples[22868]=9602;
squeal_samples[22869]=6723;
squeal_samples[22870]=5628;
squeal_samples[22871]=8487;
squeal_samples[22872]=11394;
squeal_samples[22873]=14184;
squeal_samples[22874]=16841;
squeal_samples[22875]=19395;
squeal_samples[22876]=21829;
squeal_samples[22877]=24153;
squeal_samples[22878]=26379;
squeal_samples[22879]=28501;
squeal_samples[22880]=30535;
squeal_samples[22881]=32480;
squeal_samples[22882]=34327;
squeal_samples[22883]=36105;
squeal_samples[22884]=37796;
squeal_samples[22885]=39413;
squeal_samples[22886]=40956;
squeal_samples[22887]=42429;
squeal_samples[22888]=43837;
squeal_samples[22889]=45182;
squeal_samples[22890]=46468;
squeal_samples[22891]=47697;
squeal_samples[22892]=48867;
squeal_samples[22893]=49989;
squeal_samples[22894]=51057;
squeal_samples[22895]=52081;
squeal_samples[22896]=53057;
squeal_samples[22897]=53775;
squeal_samples[22898]=49894;
squeal_samples[22899]=44417;
squeal_samples[22900]=39300;
squeal_samples[22901]=34501;
squeal_samples[22902]=30016;
squeal_samples[22903]=25818;
squeal_samples[22904]=21894;
squeal_samples[22905]=18214;
squeal_samples[22906]=14777;
squeal_samples[22907]=11550;
squeal_samples[22908]=8544;
squeal_samples[22909]=5768;
squeal_samples[22910]=6641;
squeal_samples[22911]=9623;
squeal_samples[22912]=12492;
squeal_samples[22913]=15223;
squeal_samples[22914]=17846;
squeal_samples[22915]=20345;
squeal_samples[22916]=22736;
squeal_samples[22917]=25021;
squeal_samples[22918]=27208;
squeal_samples[22919]=29297;
squeal_samples[22920]=31294;
squeal_samples[22921]=33201;
squeal_samples[22922]=35021;
squeal_samples[22923]=36766;
squeal_samples[22924]=38424;
squeal_samples[22925]=40009;
squeal_samples[22926]=41530;
squeal_samples[22927]=42977;
squeal_samples[22928]=44362;
squeal_samples[22929]=45681;
squeal_samples[22930]=46945;
squeal_samples[22931]=48151;
squeal_samples[22932]=49302;
squeal_samples[22933]=50399;
squeal_samples[22934]=51450;
squeal_samples[22935]=52454;
squeal_samples[22936]=53417;
squeal_samples[22937]=53013;
squeal_samples[22938]=47802;
squeal_samples[22939]=42454;
squeal_samples[22940]=37463;
squeal_samples[22941]=32785;
squeal_samples[22942]=28405;
squeal_samples[22943]=24312;
squeal_samples[22944]=20476;
squeal_samples[22945]=16900;
squeal_samples[22946]=13537;
squeal_samples[22947]=10401;
squeal_samples[22948]=7459;
squeal_samples[22949]=5431;
squeal_samples[22950]=7772;
squeal_samples[22951]=10710;
squeal_samples[22952]=13519;
squeal_samples[22953]=16216;
squeal_samples[22954]=18784;
squeal_samples[22955]=21250;
squeal_samples[22956]=23596;
squeal_samples[22957]=25844;
squeal_samples[22958]=27997;
squeal_samples[22959]=30047;
squeal_samples[22960]=32013;
squeal_samples[22961]=33886;
squeal_samples[22962]=35672;
squeal_samples[22963]=37390;
squeal_samples[22964]=39019;
squeal_samples[22965]=40579;
squeal_samples[22966]=42071;
squeal_samples[22967]=43491;
squeal_samples[22968]=44856;
squeal_samples[22969]=46151;
squeal_samples[22970]=47395;
squeal_samples[22971]=48580;
squeal_samples[22972]=49707;
squeal_samples[22973]=50792;
squeal_samples[22974]=51821;
squeal_samples[22975]=52809;
squeal_samples[22976]=53753;
squeal_samples[22977]=51308;
squeal_samples[22978]=45744;
squeal_samples[22979]=40535;
squeal_samples[22980]=35659;
squeal_samples[22981]=31104;
squeal_samples[22982]=26823;
squeal_samples[22983]=22834;
squeal_samples[22984]=19096;
squeal_samples[22985]=15600;
squeal_samples[22986]=12326;
squeal_samples[22987]=9263;
squeal_samples[22988]=6401;
squeal_samples[22989]=5895;
squeal_samples[22990]=8875;
squeal_samples[22991]=11769;
squeal_samples[22992]=14534;
squeal_samples[22993]=17181;
squeal_samples[22994]=19713;
squeal_samples[22995]=22134;
squeal_samples[22996]=24439;
squeal_samples[22997]=26657;
squeal_samples[22998]=28760;
squeal_samples[22999]=30785;
squeal_samples[23000]=32713;
squeal_samples[23001]=34556;
squeal_samples[23002]=36310;
squeal_samples[23003]=37996;
squeal_samples[23004]=39599;
squeal_samples[23005]=41137;
squeal_samples[23006]=42603;
squeal_samples[23007]=43999;
squeal_samples[23008]=45339;
squeal_samples[23009]=46610;
squeal_samples[23010]=47836;
squeal_samples[23011]=48995;
squeal_samples[23012]=50111;
squeal_samples[23013]=51168;
squeal_samples[23014]=52188;
squeal_samples[23015]=53156;
squeal_samples[23016]=53611;
squeal_samples[23017]=49168;
squeal_samples[23018]=43736;
squeal_samples[23019]=38660;
squeal_samples[23020]=33902;
squeal_samples[23021]=29452;
squeal_samples[23022]=25291;
squeal_samples[23023]=21395;
squeal_samples[23024]=17746;
squeal_samples[23025]=14338;
squeal_samples[23026]=11140;
squeal_samples[23027]=8156;
squeal_samples[23028]=5536;
squeal_samples[23029]=6993;
squeal_samples[23030]=9963;
squeal_samples[23031]=12806;
squeal_samples[23032]=15530;
squeal_samples[23033]=18131;
squeal_samples[23034]=20624;
squeal_samples[23035]=22991;
squeal_samples[23036]=25268;
squeal_samples[23037]=27444;
squeal_samples[23038]=29523;
squeal_samples[23039]=31502;
squeal_samples[23040]=33405;
squeal_samples[23041]=35207;
squeal_samples[23042]=36943;
squeal_samples[23043]=38594;
squeal_samples[23044]=40176;
squeal_samples[23045]=41682;
squeal_samples[23046]=43123;
squeal_samples[23047]=44493;
squeal_samples[23048]=45809;
squeal_samples[23049]=47062;
squeal_samples[23050]=48261;
squeal_samples[23051]=49410;
squeal_samples[23052]=50497;
squeal_samples[23053]=51547;
squeal_samples[23054]=52543;
squeal_samples[23055]=53500;
squeal_samples[23056]=52520;
squeal_samples[23057]=47076;
squeal_samples[23058]=41784;
squeal_samples[23059]=36826;
squeal_samples[23060]=32191;
squeal_samples[23061]=27845;
squeal_samples[23062]=23785;
squeal_samples[23063]=19987;
squeal_samples[23064]=16429;
squeal_samples[23065]=13093;
squeal_samples[23066]=9988;
squeal_samples[23067]=7068;
squeal_samples[23068]=5469;
squeal_samples[23069]=8109;
squeal_samples[23070]=11034;
squeal_samples[23071]=13832;
squeal_samples[23072]=16511;
squeal_samples[23073]=19065;
squeal_samples[23074]=21519;
squeal_samples[23075]=23846;
squeal_samples[23076]=26089;
squeal_samples[23077]=28223;
squeal_samples[23078]=30267;
squeal_samples[23079]=32211;
squeal_samples[23080]=34083;
squeal_samples[23081]=35858;
squeal_samples[23082]=37559;
squeal_samples[23083]=39187;
squeal_samples[23084]=40730;
squeal_samples[23085]=42223;
squeal_samples[23086]=43628;
squeal_samples[23087]=44985;
squeal_samples[23088]=46271;
squeal_samples[23089]=47509;
squeal_samples[23090]=48682;
squeal_samples[23091]=49811;
squeal_samples[23092]=50884;
squeal_samples[23093]=51914;
squeal_samples[23094]=52893;
squeal_samples[23095]=53782;
squeal_samples[23096]=50557;
squeal_samples[23097]=45038;
squeal_samples[23098]=39876;
squeal_samples[23099]=35038;
squeal_samples[23100]=30519;
squeal_samples[23101]=26279;
squeal_samples[23102]=22324;
squeal_samples[23103]=18612;
squeal_samples[23104]=15145;
squeal_samples[23105]=11894;
squeal_samples[23106]=8860;
squeal_samples[23107]=6014;
squeal_samples[23108]=6207;
squeal_samples[23109]=9206;
squeal_samples[23110]=12083;
squeal_samples[23111]=14835;
squeal_samples[23112]=17470;
squeal_samples[23113]=19985;
squeal_samples[23114]=22388;
squeal_samples[23115]=24685;
squeal_samples[23116]=26889;
squeal_samples[23117]=28988;
squeal_samples[23118]=30992;
squeal_samples[23119]=32913;
squeal_samples[23120]=34741;
squeal_samples[23121]=36494;
squeal_samples[23122]=38164;
squeal_samples[23123]=39763;
squeal_samples[23124]=41282;
squeal_samples[23125]=42749;
squeal_samples[23126]=44131;
squeal_samples[23127]=45467;
squeal_samples[23128]=46732;
squeal_samples[23129]=47948;
squeal_samples[23130]=49099;
squeal_samples[23131]=50213;
squeal_samples[23132]=51262;
squeal_samples[23133]=52279;
squeal_samples[23134]=53240;
squeal_samples[23135]=53321;
squeal_samples[23136]=48437;
squeal_samples[23137]=43048;
squeal_samples[23138]=38011;
squeal_samples[23139]=33296;
squeal_samples[23140]=28881;
squeal_samples[23141]=24749;
squeal_samples[23142]=20888;
squeal_samples[23143]=17271;
squeal_samples[23144]=13888;
squeal_samples[23145]=10722;
squeal_samples[23146]=7759;
squeal_samples[23147]=5394;
squeal_samples[23148]=7337;
squeal_samples[23149]=10288;
squeal_samples[23150]=13117;
squeal_samples[23151]=15825;
squeal_samples[23152]=18414;
squeal_samples[23153]=20889;
squeal_samples[23154]=23252;
squeal_samples[23155]=25513;
squeal_samples[23156]=27675;
squeal_samples[23157]=29737;
squeal_samples[23158]=31714;
squeal_samples[23159]=33593;
squeal_samples[23160]=35399;
squeal_samples[23161]=37115;
squeal_samples[23162]=38762;
squeal_samples[23163]=40330;
squeal_samples[23164]=41827;
squeal_samples[23165]=43259;
squeal_samples[23166]=44629;
squeal_samples[23167]=45933;
squeal_samples[23168]=47187;
squeal_samples[23169]=48371;
squeal_samples[23170]=49516;
squeal_samples[23171]=50598;
squeal_samples[23172]=51642;
squeal_samples[23173]=52626;
squeal_samples[23174]=53583;
squeal_samples[23175]=51915;
squeal_samples[23176]=46360;
squeal_samples[23177]=41110;
squeal_samples[23178]=36195;
squeal_samples[23179]=31596;
squeal_samples[23180]=27289;
squeal_samples[23181]=23259;
squeal_samples[23182]=19492;
squeal_samples[23183]=15968;
squeal_samples[23184]=12664;
squeal_samples[23185]=9575;
squeal_samples[23186]=6687;
squeal_samples[23187]=5589;
squeal_samples[23188]=8444;
squeal_samples[23189]=11353;
squeal_samples[23190]=14132;
squeal_samples[23191]=16802;
squeal_samples[23192]=19340;
squeal_samples[23193]=21780;
squeal_samples[23194]=24095;
squeal_samples[23195]=26324;
squeal_samples[23196]=28442;
squeal_samples[23197]=30482;
squeal_samples[23198]=32415;
squeal_samples[23199]=34274;
squeal_samples[23200]=36041;
squeal_samples[23201]=37728;
squeal_samples[23202]=39348;
squeal_samples[23203]=40886;
squeal_samples[23204]=42364;
squeal_samples[23205]=43770;
squeal_samples[23206]=45112;
squeal_samples[23207]=46399;
squeal_samples[23208]=47620;
squeal_samples[23209]=48798;
squeal_samples[23210]=49913;
squeal_samples[23211]=50981;
squeal_samples[23212]=52002;
squeal_samples[23213]=52976;
squeal_samples[23214]=53864;
squeal_samples[23215]=50625;
squeal_samples[23216]=45106;
squeal_samples[23217]=39928;
squeal_samples[23218]=35093;
squeal_samples[23219]=30562;
squeal_samples[23220]=26321;
squeal_samples[23221]=22353;
squeal_samples[23222]=18643;
squeal_samples[23223]=15167;
squeal_samples[23224]=11921;
squeal_samples[23225]=8876;
squeal_samples[23226]=6035;
squeal_samples[23227]=6219;
squeal_samples[23228]=9219;
squeal_samples[23229]=12097;
squeal_samples[23230]=14843;
squeal_samples[23231]=17474;
squeal_samples[23232]=19990;
squeal_samples[23233]=22392;
squeal_samples[23234]=24688;
squeal_samples[23235]=26884;
squeal_samples[23236]=28989;
squeal_samples[23237]=30985;
squeal_samples[23238]=32907;
squeal_samples[23239]=34737;
squeal_samples[23240]=36485;
squeal_samples[23241]=38158;
squeal_samples[23242]=39751;
squeal_samples[23243]=41278;
squeal_samples[23244]=42731;
squeal_samples[23245]=44120;
squeal_samples[23246]=45451;
squeal_samples[23247]=46715;
squeal_samples[23248]=47926;
squeal_samples[23249]=49082;
squeal_samples[23250]=50192;
squeal_samples[23251]=51244;
squeal_samples[23252]=52257;
squeal_samples[23253]=53222;
squeal_samples[23254]=53665;
squeal_samples[23255]=49215;
squeal_samples[23256]=43781;
squeal_samples[23257]=38690;
squeal_samples[23258]=33930;
squeal_samples[23259]=29475;
squeal_samples[23260]=25299;
squeal_samples[23261]=21408;
squeal_samples[23262]=17749;
squeal_samples[23263]=14334;
squeal_samples[23264]=11133;
squeal_samples[23265]=8145;
squeal_samples[23266]=5527;
squeal_samples[23267]=6973;
squeal_samples[23268]=9944;
squeal_samples[23269]=12782;
squeal_samples[23270]=15508;
squeal_samples[23271]=18105;
squeal_samples[23272]=20595;
squeal_samples[23273]=22964;
squeal_samples[23274]=25241;
squeal_samples[23275]=27411;
squeal_samples[23276]=29484;
squeal_samples[23277]=31471;
squeal_samples[23278]=33364;
squeal_samples[23279]=35172;
squeal_samples[23280]=36901;
squeal_samples[23281]=38554;
squeal_samples[23282]=40129;
squeal_samples[23283]=41642;
squeal_samples[23284]=43075;
squeal_samples[23285]=44453;
squeal_samples[23286]=45762;
squeal_samples[23287]=47020;
squeal_samples[23288]=48212;
squeal_samples[23289]=49358;
squeal_samples[23290]=50452;
squeal_samples[23291]=51493;
squeal_samples[23292]=52490;
squeal_samples[23293]=53446;
squeal_samples[23294]=53038;
squeal_samples[23295]=47813;
squeal_samples[23296]=42465;
squeal_samples[23297]=37462;
squeal_samples[23298]=32778;
squeal_samples[23299]=28392;
squeal_samples[23300]=24290;
squeal_samples[23301]=20454;
squeal_samples[23302]=16867;
squeal_samples[23303]=13503;
squeal_samples[23304]=10359;
squeal_samples[23305]=7419;
squeal_samples[23306]=5378;
squeal_samples[23307]=7720;
squeal_samples[23308]=10653;
squeal_samples[23309]=13467;
squeal_samples[23310]=16158;
squeal_samples[23311]=18728;
squeal_samples[23312]=21192;
squeal_samples[23313]=23533;
squeal_samples[23314]=25783;
squeal_samples[23315]=27925;
squeal_samples[23316]=29978;
squeal_samples[23317]=31941;
squeal_samples[23318]=33814;
squeal_samples[23319]=35600;
squeal_samples[23320]=37307;
squeal_samples[23321]=38943;
squeal_samples[23322]=40504;
squeal_samples[23323]=41991;
squeal_samples[23324]=43414;
squeal_samples[23325]=44769;
squeal_samples[23326]=46069;
squeal_samples[23327]=47308;
squeal_samples[23328]=48497;
squeal_samples[23329]=49621;
squeal_samples[23330]=50707;
squeal_samples[23331]=51732;
squeal_samples[23332]=52725;
squeal_samples[23333]=53665;
squeal_samples[23334]=51998;
squeal_samples[23335]=46429;
squeal_samples[23336]=41171;
squeal_samples[23337]=36253;
squeal_samples[23338]=31644;
squeal_samples[23339]=27329;
squeal_samples[23340]=23295;
squeal_samples[23341]=19524;
squeal_samples[23342]=15992;
squeal_samples[23343]=12682;
squeal_samples[23344]=9591;
squeal_samples[23345]=6702;
squeal_samples[23346]=5599;
squeal_samples[23347]=8453;
squeal_samples[23348]=11360;
squeal_samples[23349]=14137;
squeal_samples[23350]=16800;
squeal_samples[23351]=19339;
squeal_samples[23352]=21779;
squeal_samples[23353]=24090;
squeal_samples[23354]=26314;
squeal_samples[23355]=28435;
squeal_samples[23356]=30464;
squeal_samples[23357]=32403;
squeal_samples[23358]=34258;
squeal_samples[23359]=36025;
squeal_samples[23360]=37718;
squeal_samples[23361]=39322;
squeal_samples[23362]=40871;
squeal_samples[23363]=42340;
squeal_samples[23364]=43752;
squeal_samples[23365]=45087;
squeal_samples[23366]=46371;
squeal_samples[23367]=47598;
squeal_samples[23368]=48769;
squeal_samples[23369]=49885;
squeal_samples[23370]=50954;
squeal_samples[23371]=51971;
squeal_samples[23372]=52952;
squeal_samples[23373]=53830;
squeal_samples[23374]=50598;
squeal_samples[23375]=45071;
squeal_samples[23376]=39900;
squeal_samples[23377]=35055;
squeal_samples[23378]=30526;
squeal_samples[23379]=26285;
squeal_samples[23380]=22316;
squeal_samples[23381]=18607;
squeal_samples[23382]=15131;
squeal_samples[23383]=11879;
squeal_samples[23384]=8839;
squeal_samples[23385]=5995;
squeal_samples[23386]=6175;
squeal_samples[23387]=9179;
squeal_samples[23388]=12055;
squeal_samples[23389]=14801;
squeal_samples[23390]=17431;
squeal_samples[23391]=19950;
squeal_samples[23392]=22349;
squeal_samples[23393]=24646;
squeal_samples[23394]=26844;
squeal_samples[23395]=28945;
squeal_samples[23396]=30945;
squeal_samples[23397]=32864;
squeal_samples[23398]=34696;
squeal_samples[23399]=36444;
squeal_samples[23400]=38115;
squeal_samples[23401]=39711;
squeal_samples[23402]=41229;
squeal_samples[23403]=42690;
squeal_samples[23404]=44080;
squeal_samples[23405]=45401;
squeal_samples[23406]=46676;
squeal_samples[23407]=47882;
squeal_samples[23408]=49042;
squeal_samples[23409]=50143;
squeal_samples[23410]=51204;
squeal_samples[23411]=52209;
squeal_samples[23412]=53176;
squeal_samples[23413]=53616;
squeal_samples[23414]=49169;
squeal_samples[23415]=43733;
squeal_samples[23416]=38644;
squeal_samples[23417]=33888;
squeal_samples[23418]=29426;
squeal_samples[23419]=25260;
squeal_samples[23420]=21357;
squeal_samples[23421]=17707;
squeal_samples[23422]=14287;
squeal_samples[23423]=11091;
squeal_samples[23424]=8094;
squeal_samples[23425]=5481;
squeal_samples[23426]=6926;
squeal_samples[23427]=9897;
squeal_samples[23428]=12742;
squeal_samples[23429]=15458;
squeal_samples[23430]=18060;
squeal_samples[23431]=20547;
squeal_samples[23432]=22917;
squeal_samples[23433]=25196;
squeal_samples[23434]=27360;
squeal_samples[23435]=29447;
squeal_samples[23436]=31420;
squeal_samples[23437]=33319;
squeal_samples[23438]=35124;
squeal_samples[23439]=36854;
squeal_samples[23440]=38508;
squeal_samples[23441]=40081;
squeal_samples[23442]=41594;
squeal_samples[23443]=43030;
squeal_samples[23444]=44403;
squeal_samples[23445]=45718;
squeal_samples[23446]=46972;
squeal_samples[23447]=48163;
squeal_samples[23448]=49315;
squeal_samples[23449]=50400;
squeal_samples[23450]=51450;
squeal_samples[23451]=52441;
squeal_samples[23452]=53399;
squeal_samples[23453]=52991;
squeal_samples[23454]=47767;
squeal_samples[23455]=42415;
squeal_samples[23456]=37419;
squeal_samples[23457]=32727;
squeal_samples[23458]=28347;
squeal_samples[23459]=24242;
squeal_samples[23460]=20408;
squeal_samples[23461]=16819;
squeal_samples[23462]=13456;
squeal_samples[23463]=10312;
squeal_samples[23464]=7371;
squeal_samples[23465]=5334;
squeal_samples[23466]=7670;
squeal_samples[23467]=10606;
squeal_samples[23468]=13422;
squeal_samples[23469]=16107;
squeal_samples[23470]=18687;
squeal_samples[23471]=21139;
squeal_samples[23472]=23490;
squeal_samples[23473]=25733;
squeal_samples[23474]=27880;
squeal_samples[23475]=29930;
squeal_samples[23476]=31894;
squeal_samples[23477]=33767;
squeal_samples[23478]=35553;
squeal_samples[23479]=37260;
squeal_samples[23480]=38896;
squeal_samples[23481]=40456;
squeal_samples[23482]=41946;
squeal_samples[23483]=43365;
squeal_samples[23484]=44723;
squeal_samples[23485]=46021;
squeal_samples[23486]=47263;
squeal_samples[23487]=48447;
squeal_samples[23488]=49577;
squeal_samples[23489]=50657;
squeal_samples[23490]=51688;
squeal_samples[23491]=52674;
squeal_samples[23492]=53622;
squeal_samples[23493]=51947;
squeal_samples[23494]=46384;
squeal_samples[23495]=41125;
squeal_samples[23496]=36202;
squeal_samples[23497]=31600;
squeal_samples[23498]=27280;
squeal_samples[23499]=23249;
squeal_samples[23500]=19476;
squeal_samples[23501]=15946;
squeal_samples[23502]=12633;
squeal_samples[23503]=9547;
squeal_samples[23504]=6651;
squeal_samples[23505]=5556;
squeal_samples[23506]=8402;
squeal_samples[23507]=11315;
squeal_samples[23508]=14091;
squeal_samples[23509]=16751;
squeal_samples[23510]=19294;
squeal_samples[23511]=21728;
squeal_samples[23512]=24046;
squeal_samples[23513]=26266;
squeal_samples[23514]=28388;
squeal_samples[23515]=30418;
squeal_samples[23516]=32353;
squeal_samples[23517]=34213;
squeal_samples[23518]=35977;
squeal_samples[23519]=37671;
squeal_samples[23520]=39275;
squeal_samples[23521]=40824;
squeal_samples[23522]=42292;
squeal_samples[23523]=43704;
squeal_samples[23524]=45041;
squeal_samples[23525]=46323;
squeal_samples[23526]=47551;
squeal_samples[23527]=48721;
squeal_samples[23528]=49839;
squeal_samples[23529]=50903;
squeal_samples[23530]=51928;
squeal_samples[23531]=52900;
squeal_samples[23532]=53840;
squeal_samples[23533]=51369;
squeal_samples[23534]=45796;
squeal_samples[23535]=40575;
squeal_samples[23536]=35686;
squeal_samples[23537]=31115;
squeal_samples[23538]=26829;
squeal_samples[23539]=22822;
squeal_samples[23540]=19083;
squeal_samples[23541]=15564;
squeal_samples[23542]=12290;
squeal_samples[23543]=9215;
squeal_samples[23544]=6344;
squeal_samples[23545]=5840;
squeal_samples[23546]=8811;
squeal_samples[23547]=11697;
squeal_samples[23548]=14461;
squeal_samples[23549]=17107;
squeal_samples[23550]=19631;
squeal_samples[23551]=22048;
squeal_samples[23552]=24352;
squeal_samples[23553]=26561;
squeal_samples[23554]=28665;
squeal_samples[23555]=30692;
squeal_samples[23556]=32606;
squeal_samples[23557]=34451;
squeal_samples[23558]=36204;
squeal_samples[23559]=37890;
squeal_samples[23560]=39490;
squeal_samples[23561]=41019;
squeal_samples[23562]=42486;
squeal_samples[23563]=43877;
squeal_samples[23564]=45218;
squeal_samples[23565]=46488;
squeal_samples[23566]=47708;
squeal_samples[23567]=48867;
squeal_samples[23568]=49982;
squeal_samples[23569]=51043;
squeal_samples[23570]=52052;
squeal_samples[23571]=53024;
squeal_samples[23572]=53894;
squeal_samples[23573]=50661;
squeal_samples[23574]=45123;
squeal_samples[23575]=39946;
squeal_samples[23576]=35098;
squeal_samples[23577]=30560;
squeal_samples[23578]=26312;
squeal_samples[23579]=22339;
squeal_samples[23580]=18623;
squeal_samples[23581]=15144;
squeal_samples[23582]=11888;
squeal_samples[23583]=8842;
squeal_samples[23584]=5994;
squeal_samples[23585]=6169;
squeal_samples[23586]=9179;
squeal_samples[23587]=12038;
squeal_samples[23588]=14796;
squeal_samples[23589]=17418;
squeal_samples[23590]=19935;
squeal_samples[23591]=22328;
squeal_samples[23592]=24626;
squeal_samples[23593]=26821;
squeal_samples[23594]=28918;
squeal_samples[23595]=30927;
squeal_samples[23596]=32833;
squeal_samples[23597]=34668;
squeal_samples[23598]=36410;
squeal_samples[23599]=38083;
squeal_samples[23600]=39679;
squeal_samples[23601]=41198;
squeal_samples[23602]=42651;
squeal_samples[23603]=44043;
squeal_samples[23604]=45370;
squeal_samples[23605]=46636;
squeal_samples[23606]=47848;
squeal_samples[23607]=49001;
squeal_samples[23608]=50109;
squeal_samples[23609]=51157;
squeal_samples[23610]=52170;
squeal_samples[23611]=53128;
squeal_samples[23612]=53843;
squeal_samples[23613]=49934;
squeal_samples[23614]=44446;
squeal_samples[23615]=39312;
squeal_samples[23616]=34502;
squeal_samples[23617]=30003;
squeal_samples[23618]=25793;
squeal_samples[23619]=21851;
squeal_samples[23620]=18169;
squeal_samples[23621]=14711;
squeal_samples[23622]=11489;
squeal_samples[23623]=8463;
squeal_samples[23624]=5684;
squeal_samples[23625]=6540;
squeal_samples[23626]=9527;
squeal_samples[23627]=12385;
squeal_samples[23628]=15117;
squeal_samples[23629]=17727;
squeal_samples[23630]=20230;
squeal_samples[23631]=22606;
squeal_samples[23632]=24898;
squeal_samples[23633]=27075;
squeal_samples[23634]=29163;
squeal_samples[23635]=31156;
squeal_samples[23636]=33059;
squeal_samples[23637]=34880;
squeal_samples[23638]=36617;
squeal_samples[23639]=38273;
squeal_samples[23640]=39860;
squeal_samples[23641]=41378;
squeal_samples[23642]=42818;
squeal_samples[23643]=44200;
squeal_samples[23644]=45515;
squeal_samples[23645]=46776;
squeal_samples[23646]=47982;
squeal_samples[23647]=49132;
squeal_samples[23648]=50232;
squeal_samples[23649]=51277;
squeal_samples[23650]=52282;
squeal_samples[23651]=53236;
squeal_samples[23652]=53681;
squeal_samples[23653]=49214;
squeal_samples[23654]=43777;
squeal_samples[23655]=38683;
squeal_samples[23656]=33911;
squeal_samples[23657]=29451;
squeal_samples[23658]=25275;
squeal_samples[23659]=21366;
squeal_samples[23660]=17715;
squeal_samples[23661]=14283;
squeal_samples[23662]=11087;
squeal_samples[23663]=8088;
squeal_samples[23664]=5470;
squeal_samples[23665]=6909;
squeal_samples[23666]=9880;
squeal_samples[23667]=12720;
squeal_samples[23668]=15436;
squeal_samples[23669]=18039;
squeal_samples[23670]=20517;
squeal_samples[23671]=22892;
squeal_samples[23672]=25160;
squeal_samples[23673]=27331;
squeal_samples[23674]=29404;
squeal_samples[23675]=31386;
squeal_samples[23676]=33278;
squeal_samples[23677]=35087;
squeal_samples[23678]=36815;
squeal_samples[23679]=38469;
squeal_samples[23680]=40038;
squeal_samples[23681]=41551;
squeal_samples[23682]=42979;
squeal_samples[23683]=44357;
squeal_samples[23684]=45665;
squeal_samples[23685]=46924;
squeal_samples[23686]=48115;
squeal_samples[23687]=49257;
squeal_samples[23688]=50350;
squeal_samples[23689]=51390;
squeal_samples[23690]=52390;
squeal_samples[23691]=53340;
squeal_samples[23692]=53407;
squeal_samples[23693]=48507;
squeal_samples[23694]=43109;
squeal_samples[23695]=38056;
squeal_samples[23696]=33325;
squeal_samples[23697]=28901;
squeal_samples[23698]=24756;
squeal_samples[23699]=20887;
squeal_samples[23700]=17257;
squeal_samples[23701]=13865;
squeal_samples[23702]=10684;
squeal_samples[23703]=7721;
squeal_samples[23704]=5341;
squeal_samples[23705]=7281;
squeal_samples[23706]=10230;
squeal_samples[23707]=13058;
squeal_samples[23708]=15754;
squeal_samples[23709]=18341;
squeal_samples[23710]=20812;
squeal_samples[23711]=23166;
squeal_samples[23712]=25426;
squeal_samples[23713]=27585;
squeal_samples[23714]=29646;
squeal_samples[23715]=31621;
squeal_samples[23716]=33497;
squeal_samples[23717]=35300;
squeal_samples[23718]=37008;
squeal_samples[23719]=38658;
squeal_samples[23720]=40222;
squeal_samples[23721]=41718;
squeal_samples[23722]=43148;
squeal_samples[23723]=44510;
squeal_samples[23724]=45815;
squeal_samples[23725]=47060;
squeal_samples[23726]=48253;
squeal_samples[23727]=49385;
squeal_samples[23728]=50474;
squeal_samples[23729]=51504;
squeal_samples[23730]=52504;
squeal_samples[23731]=53441;
squeal_samples[23732]=53038;
squeal_samples[23733]=47800;
squeal_samples[23734]=42444;
squeal_samples[23735]=37437;
squeal_samples[23736]=32742;
squeal_samples[23737]=28358;
squeal_samples[23738]=24245;
squeal_samples[23739]=20407;
squeal_samples[23740]=16807;
squeal_samples[23741]=13443;
squeal_samples[23742]=10296;
squeal_samples[23743]=7347;
squeal_samples[23744]=5310;
squeal_samples[23745]=7643;
squeal_samples[23746]=10577;
squeal_samples[23747]=13388;
squeal_samples[23748]=16075;
squeal_samples[23749]=18644;
squeal_samples[23750]=21103;
squeal_samples[23751]=23443;
squeal_samples[23752]=25689;
squeal_samples[23753]=27836;
squeal_samples[23754]=29884;
squeal_samples[23755]=31846;
squeal_samples[23756]=33714;
squeal_samples[23757]=35505;
squeal_samples[23758]=37209;
squeal_samples[23759]=38846;
squeal_samples[23760]=40402;
squeal_samples[23761]=41887;
squeal_samples[23762]=43313;
squeal_samples[23763]=44665;
squeal_samples[23764]=45967;
squeal_samples[23765]=47200;
squeal_samples[23766]=48388;
squeal_samples[23767]=49514;
squeal_samples[23768]=50592;
squeal_samples[23769]=51625;
squeal_samples[23770]=52608;
squeal_samples[23771]=53555;
squeal_samples[23772]=52554;
squeal_samples[23773]=47101;
squeal_samples[23774]=41789;
squeal_samples[23775]=36825;
squeal_samples[23776]=32163;
squeal_samples[23777]=27817;
squeal_samples[23778]=23736;
squeal_samples[23779]=19936;
squeal_samples[23780]=16364;
squeal_samples[23781]=13026;
squeal_samples[23782]=9902;
squeal_samples[23783]=6984;
squeal_samples[23784]=5367;
squeal_samples[23785]=8007;
squeal_samples[23786]=10924;
squeal_samples[23787]=13718;
squeal_samples[23788]=16389;
squeal_samples[23789]=18947;
squeal_samples[23790]=21390;
squeal_samples[23791]=23719;
squeal_samples[23792]=25950;
squeal_samples[23793]=28088;
squeal_samples[23794]=30123;
squeal_samples[23795]=32072;
squeal_samples[23796]=33932;
squeal_samples[23797]=35708;
squeal_samples[23798]=37406;
squeal_samples[23799]=39027;
squeal_samples[23800]=40582;
squeal_samples[23801]=42054;
squeal_samples[23802]=43474;
squeal_samples[23803]=44817;
squeal_samples[23804]=46112;
squeal_samples[23805]=47340;
squeal_samples[23806]=48518;
squeal_samples[23807]=49638;
squeal_samples[23808]=50712;
squeal_samples[23809]=51735;
squeal_samples[23810]=52721;
squeal_samples[23811]=53652;
squeal_samples[23812]=51983;
squeal_samples[23813]=46400;
squeal_samples[23814]=41140;
squeal_samples[23815]=36211;
squeal_samples[23816]=31598;
squeal_samples[23817]=27278;
squeal_samples[23818]=23240;
squeal_samples[23819]=19460;
squeal_samples[23820]=15924;
squeal_samples[23821]=12612;
squeal_samples[23822]=9517;
squeal_samples[23823]=6615;
squeal_samples[23824]=5518;
squeal_samples[23825]=8360;
squeal_samples[23826]=11270;
squeal_samples[23827]=14046;
squeal_samples[23828]=16704;
squeal_samples[23829]=19244;
squeal_samples[23830]=21677;
squeal_samples[23831]=23995;
squeal_samples[23832]=26216;
squeal_samples[23833]=28330;
squeal_samples[23834]=30362;
squeal_samples[23835]=32298;
squeal_samples[23836]=34148;
squeal_samples[23837]=35914;
squeal_samples[23838]=37600;
squeal_samples[23839]=39216;
squeal_samples[23840]=40755;
squeal_samples[23841]=42220;
squeal_samples[23842]=43631;
squeal_samples[23843]=44975;
squeal_samples[23844]=46255;
squeal_samples[23845]=47479;
squeal_samples[23846]=48643;
squeal_samples[23847]=49763;
squeal_samples[23848]=50831;
squeal_samples[23849]=51849;
squeal_samples[23850]=52828;
squeal_samples[23851]=53757;
squeal_samples[23852]=51294;
squeal_samples[23853]=45716;
squeal_samples[23854]=40493;
squeal_samples[23855]=35601;
squeal_samples[23856]=31033;
squeal_samples[23857]=26745;
squeal_samples[23858]=22738;
squeal_samples[23859]=18994;
squeal_samples[23860]=15482;
squeal_samples[23861]=12205;
squeal_samples[23862]=9128;
squeal_samples[23863]=6258;
squeal_samples[23864]=5752;
squeal_samples[23865]=8724;
squeal_samples[23866]=11611;
squeal_samples[23867]=14374;
squeal_samples[23868]=17017;
squeal_samples[23869]=19542;
squeal_samples[23870]=21959;
squeal_samples[23871]=24264;
squeal_samples[23872]=26470;
squeal_samples[23873]=28580;
squeal_samples[23874]=30592;
squeal_samples[23875]=32523;
squeal_samples[23876]=34355;
squeal_samples[23877]=36123;
squeal_samples[23878]=37790;
squeal_samples[23879]=39402;
squeal_samples[23880]=40932;
squeal_samples[23881]=42393;
squeal_samples[23882]=43793;
squeal_samples[23883]=45125;
squeal_samples[23884]=46395;
squeal_samples[23885]=47619;
squeal_samples[23886]=48778;
squeal_samples[23887]=49887;
squeal_samples[23888]=50949;
squeal_samples[23889]=51962;
squeal_samples[23890]=52935;
squeal_samples[23891]=53854;
squeal_samples[23892]=51390;
squeal_samples[23893]=45804;
squeal_samples[23894]=40575;
squeal_samples[23895]=35680;
squeal_samples[23896]=31099;
squeal_samples[23897]=26811;
squeal_samples[23898]=22797;
squeal_samples[23899]=19051;
squeal_samples[23900]=15536;
squeal_samples[23901]=12247;
squeal_samples[23902]=9170;
squeal_samples[23903]=6297;
squeal_samples[23904]=5788;
squeal_samples[23905]=8760;
squeal_samples[23906]=11643;
squeal_samples[23907]=14405;
squeal_samples[23908]=17044;
squeal_samples[23909]=19568;
squeal_samples[23910]=21984;
squeal_samples[23911]=24287;
squeal_samples[23912]=26493;
squeal_samples[23913]=28602;
squeal_samples[23914]=30615;
squeal_samples[23915]=32538;
squeal_samples[23916]=34378;
squeal_samples[23917]=36130;
squeal_samples[23918]=37811;
squeal_samples[23919]=39411;
squeal_samples[23920]=40939;
squeal_samples[23921]=42407;
squeal_samples[23922]=43799;
squeal_samples[23923]=45137;
squeal_samples[23924]=46405;
squeal_samples[23925]=47622;
squeal_samples[23926]=48784;
squeal_samples[23927]=49890;
squeal_samples[23928]=50954;
squeal_samples[23929]=51961;
squeal_samples[23930]=52933;
squeal_samples[23931]=53860;
squeal_samples[23932]=51394;
squeal_samples[23933]=45801;
squeal_samples[23934]=40578;
squeal_samples[23935]=35679;
squeal_samples[23936]=31104;
squeal_samples[23937]=26805;
squeal_samples[23938]=22799;
squeal_samples[23939]=19043;
squeal_samples[23940]=15531;
squeal_samples[23941]=12246;
squeal_samples[23942]=9168;
squeal_samples[23943]=6292;
squeal_samples[23944]=5779;
squeal_samples[23945]=8756;
squeal_samples[23946]=11636;
squeal_samples[23947]=14399;
squeal_samples[23948]=17038;
squeal_samples[23949]=19560;
squeal_samples[23950]=21980;
squeal_samples[23951]=24278;
squeal_samples[23952]=26484;
squeal_samples[23953]=28594;
squeal_samples[23954]=30608;
squeal_samples[23955]=32529;
squeal_samples[23956]=34369;
squeal_samples[23957]=36124;
squeal_samples[23958]=37806;
squeal_samples[23959]=39401;
squeal_samples[23960]=40938;
squeal_samples[23961]=42391;
squeal_samples[23962]=43790;
squeal_samples[23963]=45122;
squeal_samples[23964]=46400;
squeal_samples[23965]=47616;
squeal_samples[23966]=48771;
squeal_samples[23967]=49887;
squeal_samples[23968]=50943;
squeal_samples[23969]=51958;
squeal_samples[23970]=52926;
squeal_samples[23971]=53846;
squeal_samples[23972]=51385;
squeal_samples[23973]=45793;
squeal_samples[23974]=40566;
squeal_samples[23975]=35670;
squeal_samples[23976]=31088;
squeal_samples[23977]=26797;
squeal_samples[23978]=22784;
squeal_samples[23979]=19034;
squeal_samples[23980]=15517;
squeal_samples[23981]=12236;
squeal_samples[23982]=9155;
squeal_samples[23983]=6285;
squeal_samples[23984]=5769;
squeal_samples[23985]=8743;
squeal_samples[23986]=11625;
squeal_samples[23987]=14387;
squeal_samples[23988]=17024;
squeal_samples[23989]=19552;
squeal_samples[23990]=21964;
squeal_samples[23991]=24269;
squeal_samples[23992]=26477;
squeal_samples[23993]=28581;
squeal_samples[23994]=30598;
squeal_samples[23995]=32515;
squeal_samples[23996]=34358;
squeal_samples[23997]=36114;
squeal_samples[23998]=37792;
squeal_samples[23999]=39391;
squeal_samples[24000]=40924;
squeal_samples[24001]=42380;
squeal_samples[24002]=43780;
squeal_samples[24003]=45108;
squeal_samples[24004]=46391;
squeal_samples[24005]=47601;
squeal_samples[24006]=48762;
squeal_samples[24007]=49873;
squeal_samples[24008]=50932;
squeal_samples[24009]=51947;
squeal_samples[24010]=52912;
squeal_samples[24011]=53837;
squeal_samples[24012]=51371;
squeal_samples[24013]=45782;
squeal_samples[24014]=40554;
squeal_samples[24015]=35658;
squeal_samples[24016]=31076;
squeal_samples[24017]=26786;
squeal_samples[24018]=22773;
squeal_samples[24019]=19024;
squeal_samples[24020]=15510;
squeal_samples[24021]=12219;
squeal_samples[24022]=9148;
squeal_samples[24023]=6271;
squeal_samples[24024]=5757;
squeal_samples[24025]=8731;
squeal_samples[24026]=11615;
squeal_samples[24027]=14372;
squeal_samples[24028]=17016;
squeal_samples[24029]=19536;
squeal_samples[24030]=21956;
squeal_samples[24031]=24255;
squeal_samples[24032]=26466;
squeal_samples[24033]=28569;
squeal_samples[24034]=30586;
squeal_samples[24035]=32510;
squeal_samples[24036]=34344;
squeal_samples[24037]=36105;
squeal_samples[24038]=37777;
squeal_samples[24039]=39384;
squeal_samples[24040]=40907;
squeal_samples[24041]=42373;
squeal_samples[24042]=43762;
squeal_samples[24043]=45104;
squeal_samples[24044]=46373;
squeal_samples[24045]=47593;
squeal_samples[24046]=48748;
squeal_samples[24047]=49861;
squeal_samples[24048]=50923;
squeal_samples[24049]=51932;
squeal_samples[24050]=52902;
squeal_samples[24051]=53825;
squeal_samples[24052]=51359;
squeal_samples[24053]=45771;
squeal_samples[24054]=40542;
squeal_samples[24055]=35645;
squeal_samples[24056]=31066;
squeal_samples[24057]=26773;
squeal_samples[24058]=22761;
squeal_samples[24059]=19014;
squeal_samples[24060]=15496;
squeal_samples[24061]=12208;
squeal_samples[24062]=9138;
squeal_samples[24063]=6255;
squeal_samples[24064]=5750;
squeal_samples[24065]=8717;
squeal_samples[24066]=11601;
squeal_samples[24067]=14366;
squeal_samples[24068]=16997;
squeal_samples[24069]=19532;
squeal_samples[24070]=21938;
squeal_samples[24071]=24247;
squeal_samples[24072]=26451;
squeal_samples[24073]=28561;
squeal_samples[24074]=30571;
squeal_samples[24075]=32501;
squeal_samples[24076]=34329;
squeal_samples[24077]=36096;
squeal_samples[24078]=37763;
squeal_samples[24079]=39374;
squeal_samples[24080]=40894;
squeal_samples[24081]=42362;
squeal_samples[24082]=43750;
squeal_samples[24083]=45091;
squeal_samples[24084]=46362;
squeal_samples[24085]=47582;
squeal_samples[24086]=48736;
squeal_samples[24087]=49849;
squeal_samples[24088]=50910;
squeal_samples[24089]=51921;
squeal_samples[24090]=52891;
squeal_samples[24091]=53813;
squeal_samples[24092]=51347;
squeal_samples[24093]=45759;
squeal_samples[24094]=40529;
squeal_samples[24095]=35637;
squeal_samples[24096]=31051;
squeal_samples[24097]=26762;
squeal_samples[24098]=22750;
squeal_samples[24099]=19001;
squeal_samples[24100]=15486;
squeal_samples[24101]=12197;
squeal_samples[24102]=9121;
squeal_samples[24103]=6250;
squeal_samples[24104]=5732;
squeal_samples[24105]=8710;
squeal_samples[24106]=11587;
squeal_samples[24107]=14354;
squeal_samples[24108]=16986;
squeal_samples[24109]=19519;
squeal_samples[24110]=21927;
squeal_samples[24111]=24236;
squeal_samples[24112]=26439;
squeal_samples[24113]=28547;
squeal_samples[24114]=30562;
squeal_samples[24115]=32486;
squeal_samples[24116]=34322;
squeal_samples[24117]=36079;
squeal_samples[24118]=37756;
squeal_samples[24119]=39357;
squeal_samples[24120]=40887;
squeal_samples[24121]=42347;
squeal_samples[24122]=43741;
squeal_samples[24123]=45078;
squeal_samples[24124]=46350;
squeal_samples[24125]=47570;
squeal_samples[24126]=48723;
squeal_samples[24127]=49840;
squeal_samples[24128]=50898;
squeal_samples[24129]=51908;
squeal_samples[24130]=52880;
squeal_samples[24131]=53799;
squeal_samples[24132]=51337;
squeal_samples[24133]=45748;
squeal_samples[24134]=40517;
squeal_samples[24135]=35624;
squeal_samples[24136]=31040;
squeal_samples[24137]=26750;
squeal_samples[24138]=22738;
squeal_samples[24139]=18990;
squeal_samples[24140]=15473;
squeal_samples[24141]=12186;
squeal_samples[24142]=9110;
squeal_samples[24143]=6237;
squeal_samples[24144]=5721;
squeal_samples[24145]=8697;
squeal_samples[24146]=11578;
squeal_samples[24147]=14339;
squeal_samples[24148]=16979;
squeal_samples[24149]=19501;
squeal_samples[24150]=21921;
squeal_samples[24151]=24219;
squeal_samples[24152]=26431;
squeal_samples[24153]=28535;
squeal_samples[24154]=30549;
squeal_samples[24155]=32475;
squeal_samples[24156]=34309;
squeal_samples[24157]=36068;
squeal_samples[24158]=37744;
squeal_samples[24159]=39346;
squeal_samples[24160]=40874;
squeal_samples[24161]=42337;
squeal_samples[24162]=43727;
squeal_samples[24163]=45068;
squeal_samples[24164]=46336;
squeal_samples[24165]=47561;
squeal_samples[24166]=48710;
squeal_samples[24167]=49828;
squeal_samples[24168]=50887;
squeal_samples[24169]=51894;
squeal_samples[24170]=52871;
squeal_samples[24171]=53786;
squeal_samples[24172]=51325;
squeal_samples[24173]=45736;
squeal_samples[24174]=40506;
squeal_samples[24175]=35611;
squeal_samples[24176]=31029;
squeal_samples[24177]=26739;
squeal_samples[24178]=22724;
squeal_samples[24179]=18980;
squeal_samples[24180]=15460;
squeal_samples[24181]=12174;
squeal_samples[24182]=9100;
squeal_samples[24183]=6223;
squeal_samples[24184]=5711;
squeal_samples[24185]=8683;
squeal_samples[24186]=11567;
squeal_samples[24187]=14327;
squeal_samples[24188]=16967;
squeal_samples[24189]=19490;
squeal_samples[24190]=21908;
squeal_samples[24191]=24208;
squeal_samples[24192]=26419;
squeal_samples[24193]=28522;
squeal_samples[24194]=30539;
squeal_samples[24195]=32462;
squeal_samples[24196]=34299;
squeal_samples[24197]=36054;
squeal_samples[24198]=37734;
squeal_samples[24199]=39332;
squeal_samples[24200]=40865;
squeal_samples[24201]=42322;
squeal_samples[24202]=43718;
squeal_samples[24203]=45053;
squeal_samples[24204]=46328;
squeal_samples[24205]=47545;
squeal_samples[24206]=48701;
squeal_samples[24207]=49814;
squeal_samples[24208]=50875;
squeal_samples[24209]=51884;
squeal_samples[24210]=52856;
squeal_samples[24211]=53775;
squeal_samples[24212]=52090;
squeal_samples[24213]=46500;
squeal_samples[24214]=41223;
squeal_samples[24215]=36277;
squeal_samples[24216]=31659;
squeal_samples[24217]=27321;
squeal_samples[24218]=23276;
squeal_samples[24219]=19486;
squeal_samples[24220]=15944;
squeal_samples[24221]=12618;
squeal_samples[24222]=9516;
squeal_samples[24223]=6609;
squeal_samples[24224]=5499;
squeal_samples[24225]=8348;
squeal_samples[24226]=11248;
squeal_samples[24227]=14020;
squeal_samples[24228]=16674;
squeal_samples[24229]=19212;
squeal_samples[24230]=21635;
squeal_samples[24231]=23952;
squeal_samples[24232]=26169;
squeal_samples[24233]=28282;
squeal_samples[24234]=30310;
squeal_samples[24235]=32244;
squeal_samples[24236]=34091;
squeal_samples[24237]=35854;
squeal_samples[24238]=37541;
squeal_samples[24239]=39149;
squeal_samples[24240]=40687;
squeal_samples[24241]=42156;
squeal_samples[24242]=43558;
squeal_samples[24243]=44899;
squeal_samples[24244]=46179;
squeal_samples[24245]=47398;
squeal_samples[24246]=48573;
squeal_samples[24247]=49681;
squeal_samples[24248]=50748;
squeal_samples[24249]=51767;
squeal_samples[24250]=52738;
squeal_samples[24251]=53665;
squeal_samples[24252]=52660;
squeal_samples[24253]=47184;
squeal_samples[24254]=41862;
squeal_samples[24255]=36882;
squeal_samples[24256]=32212;
squeal_samples[24257]=27853;
squeal_samples[24258]=23758;
squeal_samples[24259]=19947;
squeal_samples[24260]=16362;
squeal_samples[24261]=13021;
squeal_samples[24262]=9884;
squeal_samples[24263]=6957;
squeal_samples[24264]=5333;
squeal_samples[24265]=7970;
squeal_samples[24266]=10883;
squeal_samples[24267]=13677;
squeal_samples[24268]=16338;
squeal_samples[24269]=18891;
squeal_samples[24270]=21337;
squeal_samples[24271]=23657;
squeal_samples[24272]=25891;
squeal_samples[24273]=28017;
squeal_samples[24274]=30050;
squeal_samples[24275]=32001;
squeal_samples[24276]=33857;
squeal_samples[24277]=35630;
squeal_samples[24278]=37324;
squeal_samples[24279]=38947;
squeal_samples[24280]=40489;
squeal_samples[24281]=41973;
squeal_samples[24282]=43375;
squeal_samples[24283]=44729;
squeal_samples[24284]=46009;
squeal_samples[24285]=47240;
squeal_samples[24286]=48416;
squeal_samples[24287]=49536;
squeal_samples[24288]=50605;
squeal_samples[24289]=51629;
squeal_samples[24290]=52606;
squeal_samples[24291]=53546;
squeal_samples[24292]=53119;
squeal_samples[24293]=47869;
squeal_samples[24294]=42502;
squeal_samples[24295]=37476;
squeal_samples[24296]=32775;
squeal_samples[24297]=28369;
squeal_samples[24298]=24249;
squeal_samples[24299]=20399;
squeal_samples[24300]=16787;
squeal_samples[24301]=13416;
squeal_samples[24302]=10259;
squeal_samples[24303]=7301;
squeal_samples[24304]=5260;
squeal_samples[24305]=7583;
squeal_samples[24306]=10520;
squeal_samples[24307]=13316;
squeal_samples[24308]=16005;
squeal_samples[24309]=18568;
squeal_samples[24310]=21027;
squeal_samples[24311]=23364;
squeal_samples[24312]=25606;
squeal_samples[24313]=27745;
squeal_samples[24314]=29790;
squeal_samples[24315]=31751;
squeal_samples[24316]=33616;
squeal_samples[24317]=35401;
squeal_samples[24318]=37108;
squeal_samples[24319]=38730;
squeal_samples[24320]=40295;
squeal_samples[24321]=41773;
squeal_samples[24322]=43198;
squeal_samples[24323]=44549;
squeal_samples[24324]=45843;
squeal_samples[24325]=47081;
squeal_samples[24326]=48257;
squeal_samples[24327]=49388;
squeal_samples[24328]=50466;
squeal_samples[24329]=51487;
squeal_samples[24330]=52482;
squeal_samples[24331]=53412;
squeal_samples[24332]=53478;
squeal_samples[24333]=48547;
squeal_samples[24334]=43147;
squeal_samples[24335]=38069;
squeal_samples[24336]=33336;
squeal_samples[24337]=28887;
squeal_samples[24338]=24740;
squeal_samples[24339]=20851;
squeal_samples[24340]=17218;
squeal_samples[24341]=13809;
squeal_samples[24342]=10628;
squeal_samples[24343]=7650;
squeal_samples[24344]=5268;
squeal_samples[24345]=7199;
squeal_samples[24346]=10145;
squeal_samples[24347]=12967;
squeal_samples[24348]=15662;
squeal_samples[24349]=18248;
squeal_samples[24350]=20705;
squeal_samples[24351]=23069;
squeal_samples[24352]=25315;
squeal_samples[24353]=27474;
squeal_samples[24354]=29529;
squeal_samples[24355]=31498;
squeal_samples[24356]=33380;
squeal_samples[24357]=35170;
squeal_samples[24358]=36889;
squeal_samples[24359]=38522;
squeal_samples[24360]=40086;
squeal_samples[24361]=41586;
squeal_samples[24362]=43004;
squeal_samples[24363]=44375;
squeal_samples[24364]=45670;
squeal_samples[24365]=46919;
squeal_samples[24366]=48103;
squeal_samples[24367]=49237;
squeal_samples[24368]=50321;
squeal_samples[24369]=51354;
squeal_samples[24370]=52345;
squeal_samples[24371]=53291;
squeal_samples[24372]=53717;
squeal_samples[24373]=49241;
squeal_samples[24374]=43788;
squeal_samples[24375]=38675;
squeal_samples[24376]=33896;
squeal_samples[24377]=29423;
squeal_samples[24378]=25228;
squeal_samples[24379]=21318;
squeal_samples[24380]=17645;
squeal_samples[24381]=14217;
squeal_samples[24382]=10996;
squeal_samples[24383]=8001;
squeal_samples[24384]=5369;
squeal_samples[24385]=6806;
squeal_samples[24386]=9771;
squeal_samples[24387]=12605;
squeal_samples[24388]=15322;
squeal_samples[24389]=17919;
squeal_samples[24390]=20396;
squeal_samples[24391]=22763;
squeal_samples[24392]=25027;
squeal_samples[24393]=27197;
squeal_samples[24394]=29266;
squeal_samples[24395]=31246;
squeal_samples[24396]=33128;
squeal_samples[24397]=34943;
squeal_samples[24398]=36661;
squeal_samples[24399]=38311;
squeal_samples[24400]=39880;
squeal_samples[24401]=41387;
squeal_samples[24402]=42822;
squeal_samples[24403]=44192;
squeal_samples[24404]=45503;
squeal_samples[24405]=46754;
squeal_samples[24406]=47945;
squeal_samples[24407]=49092;
squeal_samples[24408]=50168;
squeal_samples[24409]=51224;
squeal_samples[24410]=52207;
squeal_samples[24411]=53165;
squeal_samples[24412]=53859;
squeal_samples[24413]=49938;
squeal_samples[24414]=44437;
squeal_samples[24415]=39284;
squeal_samples[24416]=34465;
squeal_samples[24417]=29954;
squeal_samples[24418]=25728;
squeal_samples[24419]=21782;
squeal_samples[24420]=18080;
squeal_samples[24421]=14622;
squeal_samples[24422]=11377;
squeal_samples[24423]=8353;
squeal_samples[24424]=5564;
squeal_samples[24425]=6418;
squeal_samples[24426]=9402;
squeal_samples[24427]=12244;
squeal_samples[24428]=14975;
squeal_samples[24429]=17586;
squeal_samples[24430]=20080;
squeal_samples[24431]=22465;
squeal_samples[24432]=24737;
squeal_samples[24433]=26920;
squeal_samples[24434]=28999;
squeal_samples[24435]=30994;
squeal_samples[24436]=32892;
squeal_samples[24437]=34705;
squeal_samples[24438]=36440;
squeal_samples[24439]=38097;
squeal_samples[24440]=39680;
squeal_samples[24441]=41189;
squeal_samples[24442]=42633;
squeal_samples[24443]=44010;
squeal_samples[24444]=45331;
squeal_samples[24445]=46588;
squeal_samples[24446]=47790;
squeal_samples[24447]=48933;
squeal_samples[24448]=50033;
squeal_samples[24449]=51076;
squeal_samples[24450]=52074;
squeal_samples[24451]=53038;
squeal_samples[24452]=53893;
squeal_samples[24453]=50647;
squeal_samples[24454]=45092;
squeal_samples[24455]=39902;
squeal_samples[24456]=35036;
squeal_samples[24457]=30489;
squeal_samples[24458]=26228;
squeal_samples[24459]=22241;
squeal_samples[24460]=18516;
squeal_samples[24461]=15031;
squeal_samples[24462]=11761;
squeal_samples[24463]=8706;
squeal_samples[24464]=5854;
squeal_samples[24465]=6025;
squeal_samples[24466]=9021;
squeal_samples[24467]=11884;
squeal_samples[24468]=14634;
squeal_samples[24469]=17250;
squeal_samples[24470]=19764;
squeal_samples[24471]=22156;
squeal_samples[24472]=24445;
squeal_samples[24473]=26642;
squeal_samples[24474]=28732;
squeal_samples[24475]=30739;
squeal_samples[24476]=32647;
squeal_samples[24477]=34470;
squeal_samples[24478]=36217;
squeal_samples[24479]=37885;
squeal_samples[24480]=39473;
squeal_samples[24481]=40994;
squeal_samples[24482]=42445;
squeal_samples[24483]=43833;
squeal_samples[24484]=45153;
squeal_samples[24485]=46424;
squeal_samples[24486]=47626;
squeal_samples[24487]=48786;
squeal_samples[24488]=49881;
squeal_samples[24489]=50940;
squeal_samples[24490]=51945;
squeal_samples[24491]=52903;
squeal_samples[24492]=53825;
squeal_samples[24493]=51349;
squeal_samples[24494]=45756;
squeal_samples[24495]=40520;
squeal_samples[24496]=35616;
squeal_samples[24497]=31026;
squeal_samples[24498]=26732;
squeal_samples[24499]=22712;
squeal_samples[24500]=18962;
squeal_samples[24501]=15441;
squeal_samples[24502]=12147;
squeal_samples[24503]=9063;
squeal_samples[24504]=6185;
squeal_samples[24505]=5673;
squeal_samples[24506]=8640;
squeal_samples[24507]=11525;
squeal_samples[24508]=14280;
squeal_samples[24509]=16923;
squeal_samples[24510]=19445;
squeal_samples[24511]=21857;
squeal_samples[24512]=24158;
squeal_samples[24513]=26362;
squeal_samples[24514]=28469;
squeal_samples[24515]=30474;
squeal_samples[24516]=32403;
squeal_samples[24517]=34235;
squeal_samples[24518]=35990;
squeal_samples[24519]=37665;
squeal_samples[24520]=39268;
squeal_samples[24521]=40794;
squeal_samples[24522]=42259;
squeal_samples[24523]=43648;
squeal_samples[24524]=44983;
squeal_samples[24525]=46255;
squeal_samples[24526]=47467;
squeal_samples[24527]=48629;
squeal_samples[24528]=49736;
squeal_samples[24529]=50797;
squeal_samples[24530]=51806;
squeal_samples[24531]=52778;
squeal_samples[24532]=53697;
squeal_samples[24533]=52685;
squeal_samples[24534]=47207;
squeal_samples[24535]=41875;
squeal_samples[24536]=36887;
squeal_samples[24537]=32214;
squeal_samples[24538]=27844;
squeal_samples[24539]=23755;
squeal_samples[24540]=19931;
squeal_samples[24541]=16348;
squeal_samples[24542]=12998;
squeal_samples[24543]=9862;
squeal_samples[24544]=6928;
squeal_samples[24545]=5302;
squeal_samples[24546]=7933;
squeal_samples[24547]=10850;
squeal_samples[24548]=13631;
squeal_samples[24549]=16306;
squeal_samples[24550]=18844;
squeal_samples[24551]=21294;
squeal_samples[24552]=23612;
squeal_samples[24553]=25842;
squeal_samples[24554]=27966;
squeal_samples[24555]=30004;
squeal_samples[24556]=31944;
squeal_samples[24557]=33801;
squeal_samples[24558]=35577;
squeal_samples[24559]=37269;
squeal_samples[24560]=38883;
squeal_samples[24561]=40435;
squeal_samples[24562]=41906;
squeal_samples[24563]=43319;
squeal_samples[24564]=44668;
squeal_samples[24565]=45947;
squeal_samples[24566]=47182;
squeal_samples[24567]=48348;
squeal_samples[24568]=49471;
squeal_samples[24569]=50540;
squeal_samples[24570]=51561;
squeal_samples[24571]=52542;
squeal_samples[24572]=53473;
squeal_samples[24573]=53521;
squeal_samples[24574]=48596;
squeal_samples[24575]=43180;
squeal_samples[24576]=38106;
squeal_samples[24577]=33356;
squeal_samples[24578]=28911;
squeal_samples[24579]=24747;
squeal_samples[24580]=20862;
squeal_samples[24581]=17213;
squeal_samples[24582]=13815;
squeal_samples[24583]=10619;
squeal_samples[24584]=7641;
squeal_samples[24585]=5251;
squeal_samples[24586]=7183;
squeal_samples[24587]=10124;
squeal_samples[24588]=12946;
squeal_samples[24589]=15634;
squeal_samples[24590]=18222;
squeal_samples[24591]=20677;
squeal_samples[24592]=23037;
squeal_samples[24593]=25283;
squeal_samples[24594]=27442;
squeal_samples[24595]=29496;
squeal_samples[24596]=31461;
squeal_samples[24597]=33341;
squeal_samples[24598]=35127;
squeal_samples[24599]=36848;
squeal_samples[24600]=38480;
squeal_samples[24601]=40048;
squeal_samples[24602]=41538;
squeal_samples[24603]=42959;
squeal_samples[24604]=44324;
squeal_samples[24605]=45623;
squeal_samples[24606]=46868;
squeal_samples[24607]=48053;
squeal_samples[24608]=49184;
squeal_samples[24609]=50271;
squeal_samples[24610]=51296;
squeal_samples[24611]=52293;
squeal_samples[24612]=53236;
squeal_samples[24613]=53928;
squeal_samples[24614]=49999;
squeal_samples[24615]=44485;
squeal_samples[24616]=39336;
squeal_samples[24617]=34502;
squeal_samples[24618]=29985;
squeal_samples[24619]=25749;
squeal_samples[24620]=21798;
squeal_samples[24621]=18096;
squeal_samples[24622]=14628;
squeal_samples[24623]=11391;
squeal_samples[24624]=8354;
squeal_samples[24625]=5561;
squeal_samples[24626]=6416;
squeal_samples[24627]=9388;
squeal_samples[24628]=12239;
squeal_samples[24629]=14963;
squeal_samples[24630]=17570;
squeal_samples[24631]=20069;
squeal_samples[24632]=22444;
squeal_samples[24633]=24723;
squeal_samples[24634]=26894;
squeal_samples[24635]=28983;
squeal_samples[24636]=30965;
squeal_samples[24637]=32868;
squeal_samples[24638]=34678;
squeal_samples[24639]=36415;
squeal_samples[24640]=38071;
squeal_samples[24641]=39647;
squeal_samples[24642]=41161;
squeal_samples[24643]=42598;
squeal_samples[24644]=43982;
squeal_samples[24645]=45291;
squeal_samples[24646]=46553;
squeal_samples[24647]=47752;
squeal_samples[24648]=48898;
squeal_samples[24649]=49989;
squeal_samples[24650]=51040;
squeal_samples[24651]=52037;
squeal_samples[24652]=52993;
squeal_samples[24653]=53908;
squeal_samples[24654]=51423;
squeal_samples[24655]=45816;
squeal_samples[24656]=40579;
squeal_samples[24657]=35663;
squeal_samples[24658]=31075;
squeal_samples[24659]=26770;
squeal_samples[24660]=22748;
squeal_samples[24661]=18990;
squeal_samples[24662]=15466;
squeal_samples[24663]=12169;
squeal_samples[24664]=9083;
squeal_samples[24665]=6198;
squeal_samples[24666]=5678;
squeal_samples[24667]=8647;
squeal_samples[24668]=11521;
squeal_samples[24669]=14288;
squeal_samples[24670]=16914;
squeal_samples[24671]=19447;
squeal_samples[24672]=21850;
squeal_samples[24673]=24151;
squeal_samples[24674]=26353;
squeal_samples[24675]=28453;
squeal_samples[24676]=30468;
squeal_samples[24677]=32387;
squeal_samples[24678]=34223;
squeal_samples[24679]=35974;
squeal_samples[24680]=37652;
squeal_samples[24681]=39247;
squeal_samples[24682]=40776;
squeal_samples[24683]=42238;
squeal_samples[24684]=43625;
squeal_samples[24685]=44962;
squeal_samples[24686]=46231;
squeal_samples[24687]=47441;
squeal_samples[24688]=48604;
squeal_samples[24689]=49712;
squeal_samples[24690]=50766;
squeal_samples[24691]=51778;
squeal_samples[24692]=52745;
squeal_samples[24693]=53668;
squeal_samples[24694]=52654;
squeal_samples[24695]=47177;
squeal_samples[24696]=41846;
squeal_samples[24697]=36855;
squeal_samples[24698]=32185;
squeal_samples[24699]=27807;
squeal_samples[24700]=23720;
squeal_samples[24701]=19895;
squeal_samples[24702]=16313;
squeal_samples[24703]=12962;
squeal_samples[24704]=9820;
squeal_samples[24705]=6889;
squeal_samples[24706]=5263;
squeal_samples[24707]=7896;
squeal_samples[24708]=10805;
squeal_samples[24709]=13594;
squeal_samples[24710]=16260;
squeal_samples[24711]=18812;
squeal_samples[24712]=21251;
squeal_samples[24713]=23572;
squeal_samples[24714]=25801;
squeal_samples[24715]=27924;
squeal_samples[24716]=29963;
squeal_samples[24717]=31904;
squeal_samples[24718]=33759;
squeal_samples[24719]=35537;
squeal_samples[24720]=37225;
squeal_samples[24721]=38847;
squeal_samples[24722]=40389;
squeal_samples[24723]=41868;
squeal_samples[24724]=43272;
squeal_samples[24725]=44618;
squeal_samples[24726]=45906;
squeal_samples[24727]=47131;
squeal_samples[24728]=48305;
squeal_samples[24729]=49427;
squeal_samples[24730]=50500;
squeal_samples[24731]=51521;
squeal_samples[24732]=52494;
squeal_samples[24733]=53434;
squeal_samples[24734]=53477;
squeal_samples[24735]=48553;
squeal_samples[24736]=43131;
squeal_samples[24737]=38061;
squeal_samples[24738]=33308;
squeal_samples[24739]=28865;
squeal_samples[24740]=24708;
squeal_samples[24741]=20817;
squeal_samples[24742]=17176;
squeal_samples[24743]=13765;
squeal_samples[24744]=10575;
squeal_samples[24745]=7594;
squeal_samples[24746]=5203;
squeal_samples[24747]=7140;
squeal_samples[24748]=10075;
squeal_samples[24749]=12899;
squeal_samples[24750]=15591;
squeal_samples[24751]=18171;
squeal_samples[24752]=20637;
squeal_samples[24753]=22985;
squeal_samples[24754]=25239;
squeal_samples[24755]=27395;
squeal_samples[24756]=29449;
squeal_samples[24757]=31417;
squeal_samples[24758]=33291;
squeal_samples[24759]=35084;
squeal_samples[24760]=36799;
squeal_samples[24761]=38435;
squeal_samples[24762]=40002;
squeal_samples[24763]=41489;
squeal_samples[24764]=42922;
squeal_samples[24765]=44273;
squeal_samples[24766]=45581;
squeal_samples[24767]=46819;
squeal_samples[24768]=48008;
squeal_samples[24769]=49137;
squeal_samples[24770]=50224;
squeal_samples[24771]=51256;
squeal_samples[24772]=52246;
squeal_samples[24773]=53191;
squeal_samples[24774]=53881;
squeal_samples[24775]=49951;
squeal_samples[24776]=44442;
squeal_samples[24777]=39285;
squeal_samples[24778]=34462;
squeal_samples[24779]=29932;
squeal_samples[24780]=25708;
squeal_samples[24781]=21749;
squeal_samples[24782]=18050;
squeal_samples[24783]=14584;
squeal_samples[24784]=11340;
squeal_samples[24785]=8313;
squeal_samples[24786]=5510;
squeal_samples[24787]=6373;
squeal_samples[24788]=9341;
squeal_samples[24789]=12191;
squeal_samples[24790]=14919;
squeal_samples[24791]=17522;
squeal_samples[24792]=20023;
squeal_samples[24793]=22399;
squeal_samples[24794]=24674;
squeal_samples[24795]=26850;
squeal_samples[24796]=28935;
squeal_samples[24797]=30921;
squeal_samples[24798]=32819;
squeal_samples[24799]=34634;
squeal_samples[24800]=36368;
squeal_samples[24801]=38023;
squeal_samples[24802]=39605;
squeal_samples[24803]=41109;
squeal_samples[24804]=42557;
squeal_samples[24805]=43932;
squeal_samples[24806]=45247;
squeal_samples[24807]=46505;
squeal_samples[24808]=47708;
squeal_samples[24809]=48848;
squeal_samples[24810]=49947;
squeal_samples[24811]=50989;
squeal_samples[24812]=51994;
squeal_samples[24813]=52945;
squeal_samples[24814]=53863;
squeal_samples[24815]=51374;
squeal_samples[24816]=45774;
squeal_samples[24817]=40527;
squeal_samples[24818]=35623;
squeal_samples[24819]=31024;
squeal_samples[24820]=26725;
squeal_samples[24821]=22703;
squeal_samples[24822]=18942;
squeal_samples[24823]=15421;
squeal_samples[24824]=12122;
squeal_samples[24825]=9037;
squeal_samples[24826]=6151;
squeal_samples[24827]=5633;
squeal_samples[24828]=8599;
squeal_samples[24829]=11476;
squeal_samples[24830]=14241;
squeal_samples[24831]=16869;
squeal_samples[24832]=19398;
squeal_samples[24833]=21806;
squeal_samples[24834]=24103;
squeal_samples[24835]=26308;
squeal_samples[24836]=28407;
squeal_samples[24837]=30421;
squeal_samples[24838]=32340;
squeal_samples[24839]=34178;
squeal_samples[24840]=35927;
squeal_samples[24841]=37606;
squeal_samples[24842]=39200;
squeal_samples[24843]=40731;
squeal_samples[24844]=42190;
squeal_samples[24845]=43582;
squeal_samples[24846]=44911;
squeal_samples[24847]=46188;
squeal_samples[24848]=47393;
squeal_samples[24849]=48559;
squeal_samples[24850]=49664;
squeal_samples[24851]=50720;
squeal_samples[24852]=51730;
squeal_samples[24853]=52700;
squeal_samples[24854]=53620;
squeal_samples[24855]=53183;
squeal_samples[24856]=47926;
squeal_samples[24857]=42535;
squeal_samples[24858]=37507;
squeal_samples[24859]=32782;
squeal_samples[24860]=28370;
squeal_samples[24861]=24244;
squeal_samples[24862]=20381;
squeal_samples[24863]=16766;
squeal_samples[24864]=13377;
squeal_samples[24865]=10208;
squeal_samples[24866]=7250;
squeal_samples[24867]=5197;
squeal_samples[24868]=7520;
squeal_samples[24869]=10452;
squeal_samples[24870]=13246;
squeal_samples[24871]=15929;
squeal_samples[24872]=18486;
squeal_samples[24873]=20940;
squeal_samples[24874]=23276;
squeal_samples[24875]=25514;
squeal_samples[24876]=27653;
squeal_samples[24877]=29696;
squeal_samples[24878]=31655;
squeal_samples[24879]=33509;
squeal_samples[24880]=35302;
squeal_samples[24881]=36994;
squeal_samples[24882]=38626;
squeal_samples[24883]=40177;
squeal_samples[24884]=41656;
squeal_samples[24885]=43075;
squeal_samples[24886]=44431;
squeal_samples[24887]=45722;
squeal_samples[24888]=46956;
squeal_samples[24889]=48132;
squeal_samples[24890]=49264;
squeal_samples[24891]=50336;
squeal_samples[24892]=51367;
squeal_samples[24893]=52344;
squeal_samples[24894]=53281;
squeal_samples[24895]=53973;
squeal_samples[24896]=50033;
squeal_samples[24897]=44519;
squeal_samples[24898]=39346;
squeal_samples[24899]=34519;
squeal_samples[24900]=29990;
squeal_samples[24901]=25758;
squeal_samples[24902]=21799;
squeal_samples[24903]=18089;
squeal_samples[24904]=14621;
squeal_samples[24905]=11370;
squeal_samples[24906]=8335;
squeal_samples[24907]=5534;
squeal_samples[24908]=6383;
squeal_samples[24909]=9358;
squeal_samples[24910]=12205;
squeal_samples[24911]=14930;
squeal_samples[24912]=17540;
squeal_samples[24913]=20024;
squeal_samples[24914]=22401;
squeal_samples[24915]=24681;
squeal_samples[24916]=26849;
squeal_samples[24917]=28937;
squeal_samples[24918]=30914;
squeal_samples[24919]=32822;
squeal_samples[24920]=34626;
squeal_samples[24921]=36365;
squeal_samples[24922]=38013;
squeal_samples[24923]=39597;
squeal_samples[24924]=41104;
squeal_samples[24925]=42546;
squeal_samples[24926]=43921;
squeal_samples[24927]=45233;
squeal_samples[24928]=46493;
squeal_samples[24929]=47687;
squeal_samples[24930]=48833;
squeal_samples[24931]=49930;
squeal_samples[24932]=50973;
squeal_samples[24933]=51975;
squeal_samples[24934]=52925;
squeal_samples[24935]=53839;
squeal_samples[24936]=52134;
squeal_samples[24937]=46528;
squeal_samples[24938]=41242;
squeal_samples[24939]=36279;
squeal_samples[24940]=31642;
squeal_samples[24941]=27301;
squeal_samples[24942]=23232;
squeal_samples[24943]=19446;
squeal_samples[24944]=15876;
squeal_samples[24945]=12552;
squeal_samples[24946]=9435;
squeal_samples[24947]=6524;
squeal_samples[24948]=5408;
squeal_samples[24949]=8249;
squeal_samples[24950]=11145;
squeal_samples[24951]=13908;
squeal_samples[24952]=16562;
squeal_samples[24953]=19094;
squeal_samples[24954]=21518;
squeal_samples[24955]=23825;
squeal_samples[24956]=26038;
squeal_samples[24957]=28156;
squeal_samples[24958]=30174;
squeal_samples[24959]=32106;
squeal_samples[24960]=33946;
squeal_samples[24961]=35710;
squeal_samples[24962]=37390;
squeal_samples[24963]=39000;
squeal_samples[24964]=40530;
squeal_samples[24965]=42001;
squeal_samples[24966]=43397;
squeal_samples[24967]=44739;
squeal_samples[24968]=46016;
squeal_samples[24969]=47234;
squeal_samples[24970]=48398;
squeal_samples[24971]=49513;
squeal_samples[24972]=50573;
squeal_samples[24973]=51596;
squeal_samples[24974]=52558;
squeal_samples[24975]=53494;
squeal_samples[24976]=53530;
squeal_samples[24977]=48600;
squeal_samples[24978]=43172;
squeal_samples[24979]=38090;
squeal_samples[24980]=33333;
squeal_samples[24981]=28886;
squeal_samples[24982]=24717;
squeal_samples[24983]=20826;
squeal_samples[24984]=17176;
squeal_samples[24985]=13767;
squeal_samples[24986]=10569;
squeal_samples[24987]=7586;
squeal_samples[24988]=5187;
squeal_samples[24989]=7125;
squeal_samples[24990]=10060;
squeal_samples[24991]=12879;
squeal_samples[24992]=15569;
squeal_samples[24993]=18147;
squeal_samples[24994]=20608;
squeal_samples[24995]=22963;
squeal_samples[24996]=25204;
squeal_samples[24997]=27367;
squeal_samples[24998]=29410;
squeal_samples[24999]=31382;
squeal_samples[25000]=33252;
squeal_samples[25001]=35051;
squeal_samples[25002]=36757;
squeal_samples[25003]=38398;
squeal_samples[25004]=39957;
squeal_samples[25005]=41448;
squeal_samples[25006]=42874;
squeal_samples[25007]=44231;
squeal_samples[25008]=45532;
squeal_samples[25009]=46774;
squeal_samples[25010]=47957;
squeal_samples[25011]=49093;
squeal_samples[25012]=50172;
squeal_samples[25013]=51206;
squeal_samples[25014]=52192;
squeal_samples[25015]=53136;
squeal_samples[25016]=53986;
squeal_samples[25017]=50718;
squeal_samples[25018]=45155;
squeal_samples[25019]=39945;
squeal_samples[25020]=35069;
squeal_samples[25021]=30505;
squeal_samples[25022]=26239;
squeal_samples[25023]=22242;
squeal_samples[25024]=18505;
squeal_samples[25025]=15005;
squeal_samples[25026]=11731;
squeal_samples[25027]=8672;
squeal_samples[25028]=5803;
squeal_samples[25029]=5973;
squeal_samples[25030]=8960;
squeal_samples[25031]=11821;
squeal_samples[25032]=14561;
squeal_samples[25033]=17184;
squeal_samples[25034]=19685;
squeal_samples[25035]=22076;
squeal_samples[25036]=24366;
squeal_samples[25037]=26553;
squeal_samples[25038]=28642;
squeal_samples[25039]=30641;
squeal_samples[25040]=32548;
squeal_samples[25041]=34375;
squeal_samples[25042]=36114;
squeal_samples[25043]=37781;
squeal_samples[25044]=39366;
squeal_samples[25045]=40883;
squeal_samples[25046]=42335;
squeal_samples[25047]=43716;
squeal_samples[25048]=45044;
squeal_samples[25049]=46298;
squeal_samples[25050]=47509;
squeal_samples[25051]=48660;
squeal_samples[25052]=49761;
squeal_samples[25053]=50814;
squeal_samples[25054]=51814;
squeal_samples[25055]=52778;
squeal_samples[25056]=53694;
squeal_samples[25057]=52676;
squeal_samples[25058]=47185;
squeal_samples[25059]=41847;
squeal_samples[25060]=36847;
squeal_samples[25061]=32175;
squeal_samples[25062]=27794;
squeal_samples[25063]=23699;
squeal_samples[25064]=19866;
squeal_samples[25065]=16280;
squeal_samples[25066]=12923;
squeal_samples[25067]=9781;
squeal_samples[25068]=6845;
squeal_samples[25069]=5214;
squeal_samples[25070]=7845;
squeal_samples[25071]=10751;
squeal_samples[25072]=13538;
squeal_samples[25073]=16200;
squeal_samples[25074]=18753;
squeal_samples[25075]=21183;
squeal_samples[25076]=23509;
squeal_samples[25077]=25731;
squeal_samples[25078]=27862;
squeal_samples[25079]=29889;
squeal_samples[25080]=31835;
squeal_samples[25081]=33687;
squeal_samples[25082]=35460;
squeal_samples[25083]=37148;
squeal_samples[25084]=38771;
squeal_samples[25085]=40311;
squeal_samples[25086]=41788;
squeal_samples[25087]=43194;
squeal_samples[25088]=44542;
squeal_samples[25089]=45823;
squeal_samples[25090]=47049;
squeal_samples[25091]=48222;
squeal_samples[25092]=49341;
squeal_samples[25093]=50411;
squeal_samples[25094]=51434;
squeal_samples[25095]=52405;
squeal_samples[25096]=53346;
squeal_samples[25097]=53754;
squeal_samples[25098]=49268;
squeal_samples[25099]=43796;
squeal_samples[25100]=38671;
squeal_samples[25101]=33879;
squeal_samples[25102]=29392;
squeal_samples[25103]=25188;
squeal_samples[25104]=21265;
squeal_samples[25105]=17586;
squeal_samples[25106]=14144;
squeal_samples[25107]=10925;
squeal_samples[25108]=7909;
squeal_samples[25109]=5275;
squeal_samples[25110]=6701;
squeal_samples[25111]=9669;
squeal_samples[25112]=12492;
squeal_samples[25113]=15207;
squeal_samples[25114]=17794;
squeal_samples[25115]=20273;
squeal_samples[25116]=22636;
squeal_samples[25117]=24905;
squeal_samples[25118]=27060;
squeal_samples[25119]=29131;
squeal_samples[25120]=31104;
squeal_samples[25121]=32995;
squeal_samples[25122]=34794;
squeal_samples[25123]=36516;
squeal_samples[25124]=38160;
squeal_samples[25125]=39727;
squeal_samples[25126]=41231;
squeal_samples[25127]=42663;
squeal_samples[25128]=44031;
squeal_samples[25129]=45339;
squeal_samples[25130]=46588;
squeal_samples[25131]=47775;
squeal_samples[25132]=48917;
squeal_samples[25133]=50004;
squeal_samples[25134]=51044;
squeal_samples[25135]=52039;
squeal_samples[25136]=52981;
squeal_samples[25137]=53897;
squeal_samples[25138]=51402;
squeal_samples[25139]=45793;
squeal_samples[25140]=40542;
squeal_samples[25141]=35625;
squeal_samples[25142]=31027;
squeal_samples[25143]=26717;
squeal_samples[25144]=22695;
squeal_samples[25145]=18917;
squeal_samples[25146]=15403;
squeal_samples[25147]=12093;
squeal_samples[25148]=9005;
squeal_samples[25149]=6119;
squeal_samples[25150]=5594;
squeal_samples[25151]=8562;
squeal_samples[25152]=11439;
squeal_samples[25153]=14196;
squeal_samples[25154]=16827;
squeal_samples[25155]=19350;
squeal_samples[25156]=21750;
squeal_samples[25157]=24052;
squeal_samples[25158]=26251;
squeal_samples[25159]=28354;
squeal_samples[25160]=30361;
squeal_samples[25161]=32281;
squeal_samples[25162]=34119;
squeal_samples[25163]=35866;
squeal_samples[25164]=37543;
squeal_samples[25165]=39134;
squeal_samples[25166]=40666;
squeal_samples[25167]=42121;
squeal_samples[25168]=43513;
squeal_samples[25169]=44847;
squeal_samples[25170]=46111;
squeal_samples[25171]=47329;
squeal_samples[25172]=48483;
squeal_samples[25173]=49593;
squeal_samples[25174]=50646;
squeal_samples[25175]=51662;
squeal_samples[25176]=52623;
squeal_samples[25177]=53545;
squeal_samples[25178]=53108;
squeal_samples[25179]=47842;
squeal_samples[25180]=42457;
squeal_samples[25181]=37423;
squeal_samples[25182]=32703;
squeal_samples[25183]=28289;
squeal_samples[25184]=24161;
squeal_samples[25185]=20296;
squeal_samples[25186]=16679;
squeal_samples[25187]=13294;
squeal_samples[25188]=10131;
squeal_samples[25189]=7164;
squeal_samples[25190]=5114;
squeal_samples[25191]=7433;
squeal_samples[25192]=10364;
squeal_samples[25193]=13162;
squeal_samples[25194]=15838;
squeal_samples[25195]=18404;
squeal_samples[25196]=20851;
squeal_samples[25197]=23191;
squeal_samples[25198]=25426;
squeal_samples[25199]=27567;
squeal_samples[25200]=29609;
squeal_samples[25201]=31564;
squeal_samples[25202]=33422;
squeal_samples[25203]=35210;
squeal_samples[25204]=36907;
squeal_samples[25205]=38541;
squeal_samples[25206]=40088;
squeal_samples[25207]=41572;
squeal_samples[25208]=42988;
squeal_samples[25209]=44337;
squeal_samples[25210]=45634;
squeal_samples[25211]=46865;
squeal_samples[25212]=48049;
squeal_samples[25213]=49168;
squeal_samples[25214]=50247;
squeal_samples[25215]=51274;
squeal_samples[25216]=52250;
squeal_samples[25217]=53198;
squeal_samples[25218]=54030;
squeal_samples[25219]=50771;
squeal_samples[25220]=45189;
squeal_samples[25221]=39984;
squeal_samples[25222]=35095;
squeal_samples[25223]=30532;
squeal_samples[25224]=26250;
squeal_samples[25225]=22250;
squeal_samples[25226]=18513;
squeal_samples[25227]=15012;
squeal_samples[25228]=11730;
squeal_samples[25229]=8667;
squeal_samples[25230]=5795;
squeal_samples[25231]=5958;
squeal_samples[25232]=8952;
squeal_samples[25233]=11806;
squeal_samples[25234]=14550;
squeal_samples[25235]=17160;
squeal_samples[25236]=19669;
squeal_samples[25237]=22054;
squeal_samples[25238]=24342;
squeal_samples[25239]=26527;
squeal_samples[25240]=28619;
squeal_samples[25241]=30613;
squeal_samples[25242]=32522;
squeal_samples[25243]=34340;
squeal_samples[25244]=36087;
squeal_samples[25245]=37743;
squeal_samples[25246]=39337;
squeal_samples[25247]=40847;
squeal_samples[25248]=42299;
squeal_samples[25249]=43681;
squeal_samples[25250]=45000;
squeal_samples[25251]=46265;
squeal_samples[25252]=47470;
squeal_samples[25253]=48622;
squeal_samples[25254]=49717;
squeal_samples[25255]=50768;
squeal_samples[25256]=51772;
squeal_samples[25257]=52731;
squeal_samples[25258]=53646;
squeal_samples[25259]=53205;
squeal_samples[25260]=47932;
squeal_samples[25261]=42544;
squeal_samples[25262]=37496;
squeal_samples[25263]=32773;
squeal_samples[25264]=28352;
squeal_samples[25265]=24215;
squeal_samples[25266]=20347;
squeal_samples[25267]=16729;
squeal_samples[25268]=13334;
squeal_samples[25269]=10168;
squeal_samples[25270]=7196;
squeal_samples[25271]=5144;
squeal_samples[25272]=7464;
squeal_samples[25273]=10391;
squeal_samples[25274]=13186;
squeal_samples[25275]=15866;
squeal_samples[25276]=18423;
squeal_samples[25277]=20871;
squeal_samples[25278]=23206;
squeal_samples[25279]=25442;
squeal_samples[25280]=27581;
squeal_samples[25281]=29621;
squeal_samples[25282]=31569;
squeal_samples[25283]=33436;
squeal_samples[25284]=35216;
squeal_samples[25285]=36914;
squeal_samples[25286]=38543;
squeal_samples[25287]=40092;
squeal_samples[25288]=41578;
squeal_samples[25289]=42984;
squeal_samples[25290]=44344;
squeal_samples[25291]=45630;
squeal_samples[25292]=46864;
squeal_samples[25293]=48044;
squeal_samples[25294]=49164;
squeal_samples[25295]=50243;
squeal_samples[25296]=51265;
squeal_samples[25297]=52245;
squeal_samples[25298]=53190;
squeal_samples[25299]=54024;
squeal_samples[25300]=50758;
squeal_samples[25301]=45179;
squeal_samples[25302]=39970;
squeal_samples[25303]=35083;
squeal_samples[25304]=30521;
squeal_samples[25305]=26236;
squeal_samples[25306]=22241;
squeal_samples[25307]=18493;
squeal_samples[25308]=14994;
squeal_samples[25309]=11714;
squeal_samples[25310]=8647;
squeal_samples[25311]=5780;
squeal_samples[25312]=5939;
squeal_samples[25313]=8935;
squeal_samples[25314]=11789;
squeal_samples[25315]=14529;
squeal_samples[25316]=17147;
squeal_samples[25317]=19648;
squeal_samples[25318]=22039;
squeal_samples[25319]=24323;
squeal_samples[25320]=26510;
squeal_samples[25321]=28602;
squeal_samples[25322]=30595;
squeal_samples[25323]=32504;
squeal_samples[25324]=34323;
squeal_samples[25325]=36064;
squeal_samples[25326]=37726;
squeal_samples[25327]=39312;
squeal_samples[25328]=40832;
squeal_samples[25329]=42278;
squeal_samples[25330]=43662;
squeal_samples[25331]=44980;
squeal_samples[25332]=46243;
squeal_samples[25333]=47447;
squeal_samples[25334]=48598;
squeal_samples[25335]=49701;
squeal_samples[25336]=50750;
squeal_samples[25337]=51749;
squeal_samples[25338]=52714;
squeal_samples[25339]=53628;
squeal_samples[25340]=53182;
squeal_samples[25341]=47909;
squeal_samples[25342]=42521;
squeal_samples[25343]=37473;
squeal_samples[25344]=32756;
squeal_samples[25345]=28333;
squeal_samples[25346]=24198;
squeal_samples[25347]=20330;
squeal_samples[25348]=16704;
squeal_samples[25349]=13314;
squeal_samples[25350]=10143;
squeal_samples[25351]=7179;
squeal_samples[25352]=5121;
squeal_samples[25353]=7441;
squeal_samples[25354]=10367;
squeal_samples[25355]=13165;
squeal_samples[25356]=15842;
squeal_samples[25357]=18400;
squeal_samples[25358]=20848;
squeal_samples[25359]=23183;
squeal_samples[25360]=25419;
squeal_samples[25361]=27558;
squeal_samples[25362]=29597;
squeal_samples[25363]=31548;
squeal_samples[25364]=33411;
squeal_samples[25365]=35195;
squeal_samples[25366]=36889;
squeal_samples[25367]=38520;
squeal_samples[25368]=40070;
squeal_samples[25369]=41554;
squeal_samples[25370]=42967;
squeal_samples[25371]=44321;
squeal_samples[25372]=45605;
squeal_samples[25373]=46845;
squeal_samples[25374]=48016;
squeal_samples[25375]=49146;
squeal_samples[25376]=50217;
squeal_samples[25377]=51242;
squeal_samples[25378]=52229;
squeal_samples[25379]=53164;
squeal_samples[25380]=54006;
squeal_samples[25381]=50729;
squeal_samples[25382]=45161;
squeal_samples[25383]=39943;
squeal_samples[25384]=35064;
squeal_samples[25385]=30493;
squeal_samples[25386]=26217;
squeal_samples[25387]=22215;
squeal_samples[25388]=18472;
squeal_samples[25389]=14971;
squeal_samples[25390]=11690;
squeal_samples[25391]=8624;
squeal_samples[25392]=5758;
squeal_samples[25393]=5915;
squeal_samples[25394]=8913;
squeal_samples[25395]=11764;
squeal_samples[25396]=14510;
squeal_samples[25397]=17119;
squeal_samples[25398]=19630;
squeal_samples[25399]=22011;
squeal_samples[25400]=24304;
squeal_samples[25401]=26485;
squeal_samples[25402]=28579;
squeal_samples[25403]=30573;
squeal_samples[25404]=32479;
squeal_samples[25405]=34303;
squeal_samples[25406]=36038;
squeal_samples[25407]=37705;
squeal_samples[25408]=39288;
squeal_samples[25409]=40810;
squeal_samples[25410]=42255;
squeal_samples[25411]=43643;
squeal_samples[25412]=44958;
squeal_samples[25413]=46220;
squeal_samples[25414]=47424;
squeal_samples[25415]=48575;
squeal_samples[25416]=49678;
squeal_samples[25417]=50726;
squeal_samples[25418]=51726;
squeal_samples[25419]=52692;
squeal_samples[25420]=53604;
squeal_samples[25421]=53160;
squeal_samples[25422]=47886;
squeal_samples[25423]=42496;
squeal_samples[25424]=37453;
squeal_samples[25425]=32730;
squeal_samples[25426]=28313;
squeal_samples[25427]=24173;
squeal_samples[25428]=20307;
squeal_samples[25429]=16683;
squeal_samples[25430]=13288;
squeal_samples[25431]=10122;
squeal_samples[25432]=7156;
squeal_samples[25433]=5096;
squeal_samples[25434]=7420;
squeal_samples[25435]=10344;
squeal_samples[25436]=13140;
squeal_samples[25437]=15821;
squeal_samples[25438]=18376;
squeal_samples[25439]=20824;
squeal_samples[25440]=23163;
squeal_samples[25441]=25393;
squeal_samples[25442]=27536;
squeal_samples[25443]=29575;
squeal_samples[25444]=31522;
squeal_samples[25445]=33391;
squeal_samples[25446]=35170;
squeal_samples[25447]=36867;
squeal_samples[25448]=38498;
squeal_samples[25449]=40045;
squeal_samples[25450]=41532;
squeal_samples[25451]=42944;
squeal_samples[25452]=44298;
squeal_samples[25453]=45583;
squeal_samples[25454]=46820;
squeal_samples[25455]=47994;
squeal_samples[25456]=49124;
squeal_samples[25457]=50191;
squeal_samples[25458]=51224;
squeal_samples[25459]=52201;
squeal_samples[25460]=53144;
squeal_samples[25461]=53982;
squeal_samples[25462]=50706;
squeal_samples[25463]=45138;
squeal_samples[25464]=39920;
squeal_samples[25465]=35041;
squeal_samples[25466]=30470;
squeal_samples[25467]=26196;
squeal_samples[25468]=22188;
squeal_samples[25469]=18453;
squeal_samples[25470]=14945;
squeal_samples[25471]=11668;
squeal_samples[25472]=8603;
squeal_samples[25473]=5730;
squeal_samples[25474]=5899;
squeal_samples[25475]=8882;
squeal_samples[25476]=11749;
squeal_samples[25477]=14480;
squeal_samples[25478]=17101;
squeal_samples[25479]=19603;
squeal_samples[25480]=21991;
squeal_samples[25481]=24279;
squeal_samples[25482]=26463;
squeal_samples[25483]=28556;
squeal_samples[25484]=30549;
squeal_samples[25485]=32457;
squeal_samples[25486]=34279;
squeal_samples[25487]=36015;
squeal_samples[25488]=37683;
squeal_samples[25489]=39264;
squeal_samples[25490]=40787;
squeal_samples[25491]=42233;
squeal_samples[25492]=43618;
squeal_samples[25493]=44937;
squeal_samples[25494]=46196;
squeal_samples[25495]=47400;
squeal_samples[25496]=48554;
squeal_samples[25497]=49652;
squeal_samples[25498]=50706;
squeal_samples[25499]=51702;
squeal_samples[25500]=52667;
squeal_samples[25501]=53584;
squeal_samples[25502]=53134;
squeal_samples[25503]=47865;
squeal_samples[25504]=42473;
squeal_samples[25505]=37429;
squeal_samples[25506]=32707;
squeal_samples[25507]=28291;
squeal_samples[25508]=24148;
squeal_samples[25509]=20288;
squeal_samples[25510]=16654;
squeal_samples[25511]=13271;
squeal_samples[25512]=10095;
squeal_samples[25513]=7134;
squeal_samples[25514]=5074;
squeal_samples[25515]=7394;
squeal_samples[25516]=10324;
squeal_samples[25517]=13116;
squeal_samples[25518]=15797;
squeal_samples[25519]=18354;
squeal_samples[25520]=20800;
squeal_samples[25521]=23140;
squeal_samples[25522]=25370;
squeal_samples[25523]=27514;
squeal_samples[25524]=29550;
squeal_samples[25525]=31500;
squeal_samples[25526]=33369;
squeal_samples[25527]=35143;
squeal_samples[25528]=36849;
squeal_samples[25529]=38469;
squeal_samples[25530]=40028;
squeal_samples[25531]=41504;
squeal_samples[25532]=42923;
squeal_samples[25533]=44275;
squeal_samples[25534]=45557;
squeal_samples[25535]=46801;
squeal_samples[25536]=47967;
squeal_samples[25537]=49102;
squeal_samples[25538]=50169;
squeal_samples[25539]=51197;
squeal_samples[25540]=52182;
squeal_samples[25541]=53117;
squeal_samples[25542]=54014;
squeal_samples[25543]=51508;
squeal_samples[25544]=45886;
squeal_samples[25545]=40620;
squeal_samples[25546]=35696;
squeal_samples[25547]=31082;
squeal_samples[25548]=26769;
squeal_samples[25549]=22725;
squeal_samples[25550]=18951;
squeal_samples[25551]=15409;
squeal_samples[25552]=12104;
squeal_samples[25553]=8999;
squeal_samples[25554]=6109;
squeal_samples[25555]=5582;
squeal_samples[25556]=8543;
squeal_samples[25557]=11417;
squeal_samples[25558]=14167;
squeal_samples[25559]=16793;
squeal_samples[25560]=19316;
squeal_samples[25561]=21711;
squeal_samples[25562]=24012;
squeal_samples[25563]=26206;
squeal_samples[25564]=28310;
squeal_samples[25565]=30310;
squeal_samples[25566]=32226;
squeal_samples[25567]=34062;
squeal_samples[25568]=35805;
squeal_samples[25569]=37482;
squeal_samples[25570]=39073;
squeal_samples[25571]=40599;
squeal_samples[25572]=42054;
squeal_samples[25573]=43442;
squeal_samples[25574]=44772;
squeal_samples[25575]=46038;
squeal_samples[25576]=47247;
squeal_samples[25577]=48403;
squeal_samples[25578]=49513;
squeal_samples[25579]=50564;
squeal_samples[25580]=51578;
squeal_samples[25581]=52539;
squeal_samples[25582]=53461;
squeal_samples[25583]=53862;
squeal_samples[25584]=49354;
squeal_samples[25585]=43878;
squeal_samples[25586]=38729;
squeal_samples[25587]=33935;
squeal_samples[25588]=29423;
squeal_samples[25589]=25215;
squeal_samples[25590]=21278;
squeal_samples[25591]=17586;
squeal_samples[25592]=14145;
squeal_samples[25593]=10907;
squeal_samples[25594]=7889;
squeal_samples[25595]=5246;
squeal_samples[25596]=6675;
squeal_samples[25597]=9631;
squeal_samples[25598]=12453;
squeal_samples[25599]=15159;
squeal_samples[25600]=17744;
squeal_samples[25601]=20220;
squeal_samples[25602]=22575;
squeal_samples[25603]=24841;
squeal_samples[25604]=26998;
squeal_samples[25605]=29064;
squeal_samples[25606]=31029;
squeal_samples[25607]=32917;
squeal_samples[25608]=34714;
squeal_samples[25609]=36439;
squeal_samples[25610]=38074;
squeal_samples[25611]=39644;
squeal_samples[25612]=41140;
squeal_samples[25613]=42574;
squeal_samples[25614]=43941;
squeal_samples[25615]=45243;
squeal_samples[25616]=46494;
squeal_samples[25617]=47679;
squeal_samples[25618]=48817;
squeal_samples[25619]=49901;
squeal_samples[25620]=50940;
squeal_samples[25621]=51930;
squeal_samples[25622]=52877;
squeal_samples[25623]=53781;
squeal_samples[25624]=52754;
squeal_samples[25625]=47245;
squeal_samples[25626]=41897;
squeal_samples[25627]=36883;
squeal_samples[25628]=32194;
squeal_samples[25629]=27805;
squeal_samples[25630]=23695;
squeal_samples[25631]=19862;
squeal_samples[25632]=16255;
squeal_samples[25633]=12895;
squeal_samples[25634]=9742;
squeal_samples[25635]=6799;
squeal_samples[25636]=5159;
squeal_samples[25637]=7789;
squeal_samples[25638]=10691;
squeal_samples[25639]=13475;
squeal_samples[25640]=16131;
squeal_samples[25641]=18676;
squeal_samples[25642]=21111;
squeal_samples[25643]=23427;
squeal_samples[25644]=25646;
squeal_samples[25645]=27771;
squeal_samples[25646]=29797;
squeal_samples[25647]=31740;
squeal_samples[25648]=33589;
squeal_samples[25649]=35365;
squeal_samples[25650]=37044;
squeal_samples[25651]=38665;
squeal_samples[25652]=40198;
squeal_samples[25653]=41680;
squeal_samples[25654]=43081;
squeal_samples[25655]=44425;
squeal_samples[25656]=45702;
squeal_samples[25657]=46934;
squeal_samples[25658]=48100;
squeal_samples[25659]=49220;
squeal_samples[25660]=50285;
squeal_samples[25661]=51305;
squeal_samples[25662]=52281;
squeal_samples[25663]=53214;
squeal_samples[25664]=54050;
squeal_samples[25665]=50767;
squeal_samples[25666]=45189;
squeal_samples[25667]=39965;
squeal_samples[25668]=35078;
squeal_samples[25669]=30504;
squeal_samples[25670]=26217;
squeal_samples[25671]=22220;
squeal_samples[25672]=18464;
squeal_samples[25673]=14961;
squeal_samples[25674]=11674;
squeal_samples[25675]=8604;
squeal_samples[25676]=5728;
squeal_samples[25677]=5892;
squeal_samples[25678]=8877;
squeal_samples[25679]=11735;
squeal_samples[25680]=14475;
squeal_samples[25681]=17084;
squeal_samples[25682]=19589;
squeal_samples[25683]=21977;
squeal_samples[25684]=24264;
squeal_samples[25685]=26442;
squeal_samples[25686]=28536;
squeal_samples[25687]=30525;
squeal_samples[25688]=32430;
squeal_samples[25689]=34255;
squeal_samples[25690]=35989;
squeal_samples[25691]=37651;
squeal_samples[25692]=39235;
squeal_samples[25693]=40753;
squeal_samples[25694]=42200;
squeal_samples[25695]=43578;
squeal_samples[25696]=44905;
squeal_samples[25697]=46155;
squeal_samples[25698]=47367;
squeal_samples[25699]=48515;
squeal_samples[25700]=49611;
squeal_samples[25701]=50665;
squeal_samples[25702]=51662;
squeal_samples[25703]=52630;
squeal_samples[25704]=53536;
squeal_samples[25705]=53569;
squeal_samples[25706]=48620;
squeal_samples[25707]=43175;
squeal_samples[25708]=38083;
squeal_samples[25709]=33312;
squeal_samples[25710]=28854;
squeal_samples[25711]=24676;
squeal_samples[25712]=20767;
squeal_samples[25713]=17116;
squeal_samples[25714]=13688;
squeal_samples[25715]=10488;
squeal_samples[25716]=7496;
squeal_samples[25717]=5096;
squeal_samples[25718]=7016;
squeal_samples[25719]=9954;
squeal_samples[25720]=12766;
squeal_samples[25721]=15456;
squeal_samples[25722]=18030;
squeal_samples[25723]=20488;
squeal_samples[25724]=22835;
squeal_samples[25725]=25081;
squeal_samples[25726]=27226;
squeal_samples[25727]=29276;
squeal_samples[25728]=31242;
squeal_samples[25729]=33113;
squeal_samples[25730]=34897;
squeal_samples[25731]=36611;
squeal_samples[25732]=38238;
squeal_samples[25733]=39807;
squeal_samples[25734]=41288;
squeal_samples[25735]=42714;
squeal_samples[25736]=44067;
squeal_samples[25737]=45369;
squeal_samples[25738]=46607;
squeal_samples[25739]=47794;
squeal_samples[25740]=48921;
squeal_samples[25741]=50003;
squeal_samples[25742]=51031;
squeal_samples[25743]=52019;
squeal_samples[25744]=52962;
squeal_samples[25745]=53861;
squeal_samples[25746]=52143;
squeal_samples[25747]=46526;
squeal_samples[25748]=41216;
squeal_samples[25749]=36244;
squeal_samples[25750]=31595;
squeal_samples[25751]=27244;
squeal_samples[25752]=23166;
squeal_samples[25753]=19358;
squeal_samples[25754]=15790;
squeal_samples[25755]=12453;
squeal_samples[25756]=9332;
squeal_samples[25757]=6407;
squeal_samples[25758]=5284;
squeal_samples[25759]=8122;
squeal_samples[25760]=11011;
squeal_samples[25761]=13776;
squeal_samples[25762]=16423;
squeal_samples[25763]=18950;
squeal_samples[25764]=21369;
squeal_samples[25765]=23674;
squeal_samples[25766]=25884;
squeal_samples[25767]=27995;
squeal_samples[25768]=30014;
squeal_samples[25769]=31941;
squeal_samples[25770]=33780;
squeal_samples[25771]=35537;
squeal_samples[25772]=37221;
squeal_samples[25773]=38826;
squeal_samples[25774]=40356;
squeal_samples[25775]=41824;
squeal_samples[25776]=43213;
squeal_samples[25777]=44554;
squeal_samples[25778]=45825;
squeal_samples[25779]=47049;
squeal_samples[25780]=48209;
squeal_samples[25781]=49320;
squeal_samples[25782]=50379;
squeal_samples[25783]=51398;
squeal_samples[25784]=52357;
squeal_samples[25785]=53293;
squeal_samples[25786]=53961;
squeal_samples[25787]=50019;
squeal_samples[25788]=44483;
squeal_samples[25789]=39301;
squeal_samples[25790]=34460;
squeal_samples[25791]=29914;
squeal_samples[25792]=25673;
squeal_samples[25793]=21696;
squeal_samples[25794]=17982;
squeal_samples[25795]=14503;
squeal_samples[25796]=11246;
squeal_samples[25797]=8201;
squeal_samples[25798]=5392;
squeal_samples[25799]=6240;
squeal_samples[25800]=9205;
squeal_samples[25801]=12049;
squeal_samples[25802]=14770;
squeal_samples[25803]=17370;
squeal_samples[25804]=19859;
squeal_samples[25805]=22229;
squeal_samples[25806]=24505;
squeal_samples[25807]=26675;
squeal_samples[25808]=28749;
squeal_samples[25809]=30736;
squeal_samples[25810]=32627;
squeal_samples[25811]=34437;
squeal_samples[25812]=36166;
squeal_samples[25813]=37816;
squeal_samples[25814]=39397;
squeal_samples[25815]=40901;
squeal_samples[25816]=42344;
squeal_samples[25817]=43713;
squeal_samples[25818]=45030;
squeal_samples[25819]=46280;
squeal_samples[25820]=47478;
squeal_samples[25821]=48619;
squeal_samples[25822]=49717;
squeal_samples[25823]=50755;
squeal_samples[25824]=51752;
squeal_samples[25825]=52704;
squeal_samples[25826]=53614;
squeal_samples[25827]=53168;
squeal_samples[25828]=47885;
squeal_samples[25829]=42488;
squeal_samples[25830]=37434;
squeal_samples[25831]=32707;
squeal_samples[25832]=28281;
squeal_samples[25833]=24141;
squeal_samples[25834]=20266;
squeal_samples[25835]=16641;
squeal_samples[25836]=13247;
squeal_samples[25837]=10066;
squeal_samples[25838]=7096;
squeal_samples[25839]=5035;
squeal_samples[25840]=7356;
squeal_samples[25841]=10278;
squeal_samples[25842]=13073;
squeal_samples[25843]=15747;
squeal_samples[25844]=18303;
squeal_samples[25845]=20754;
squeal_samples[25846]=23080;
squeal_samples[25847]=25318;
squeal_samples[25848]=27452;
squeal_samples[25849]=29489;
squeal_samples[25850]=31448;
squeal_samples[25851]=33303;
squeal_samples[25852]=35089;
squeal_samples[25853]=36782;
squeal_samples[25854]=38408;
squeal_samples[25855]=39958;
squeal_samples[25856]=41435;
squeal_samples[25857]=42852;
squeal_samples[25858]=44201;
squeal_samples[25859]=45494;
squeal_samples[25860]=46721;
squeal_samples[25861]=47898;
squeal_samples[25862]=49022;
squeal_samples[25863]=50101;
squeal_samples[25864]=51116;
squeal_samples[25865]=52108;
squeal_samples[25866]=53036;
squeal_samples[25867]=53939;
squeal_samples[25868]=52207;
squeal_samples[25869]=46587;
squeal_samples[25870]=41269;
squeal_samples[25871]=36299;
squeal_samples[25872]=31634;
squeal_samples[25873]=27286;
squeal_samples[25874]=23194;
squeal_samples[25875]=19391;
squeal_samples[25876]=15817;
squeal_samples[25877]=12473;
squeal_samples[25878]=9352;
squeal_samples[25879]=6418;
squeal_samples[25880]=5296;
squeal_samples[25881]=8134;
squeal_samples[25882]=11017;
squeal_samples[25883]=13789;
squeal_samples[25884]=16421;
squeal_samples[25885]=18956;
squeal_samples[25886]=21371;
squeal_samples[25887]=23669;
squeal_samples[25888]=25887;
squeal_samples[25889]=27987;
squeal_samples[25890]=30010;
squeal_samples[25891]=31929;
squeal_samples[25892]=33774;
squeal_samples[25893]=35529;
squeal_samples[25894]=37208;
squeal_samples[25895]=38812;
squeal_samples[25896]=40343;
squeal_samples[25897]=41809;
squeal_samples[25898]=43201;
squeal_samples[25899]=44539;
squeal_samples[25900]=45813;
squeal_samples[25901]=47029;
squeal_samples[25902]=48191;
squeal_samples[25903]=49299;
squeal_samples[25904]=50362;
squeal_samples[25905]=51376;
squeal_samples[25906]=52341;
squeal_samples[25907]=53270;
squeal_samples[25908]=54097;
squeal_samples[25909]=50814;
squeal_samples[25910]=45223;
squeal_samples[25911]=39996;
squeal_samples[25912]=35100;
squeal_samples[25913]=30524;
squeal_samples[25914]=26231;
squeal_samples[25915]=22224;
squeal_samples[25916]=18464;
squeal_samples[25917]=14959;
squeal_samples[25918]=11666;
squeal_samples[25919]=8595;
squeal_samples[25920]=5718;
squeal_samples[25921]=5874;
squeal_samples[25922]=8864;
squeal_samples[25923]=11711;
squeal_samples[25924]=14450;
squeal_samples[25925]=17056;
squeal_samples[25926]=19563;
squeal_samples[25927]=21946;
squeal_samples[25928]=24228;
squeal_samples[25929]=26414;
squeal_samples[25930]=28495;
squeal_samples[25931]=30489;
squeal_samples[25932]=32393;
squeal_samples[25933]=34210;
squeal_samples[25934]=35946;
squeal_samples[25935]=37609;
squeal_samples[25936]=39190;
squeal_samples[25937]=40707;
squeal_samples[25938]=42154;
squeal_samples[25939]=43533;
squeal_samples[25940]=44852;
squeal_samples[25941]=46110;
squeal_samples[25942]=47316;
squeal_samples[25943]=48462;
squeal_samples[25944]=49558;
squeal_samples[25945]=50609;
squeal_samples[25946]=51610;
squeal_samples[25947]=52573;
squeal_samples[25948]=53483;
squeal_samples[25949]=53883;
squeal_samples[25950]=49371;
squeal_samples[25951]=43876;
squeal_samples[25952]=38734;
squeal_samples[25953]=33915;
squeal_samples[25954]=29411;
squeal_samples[25955]=25193;
squeal_samples[25956]=21255;
squeal_samples[25957]=17558;
squeal_samples[25958]=14104;
squeal_samples[25959]=10868;
squeal_samples[25960]=7844;
squeal_samples[25961]=5193;
squeal_samples[25962]=6621;
squeal_samples[25963]=9573;
squeal_samples[25964]=12397;
squeal_samples[25965]=15104;
squeal_samples[25966]=17686;
squeal_samples[25967]=20159;
squeal_samples[25968]=22514;
squeal_samples[25969]=24773;
squeal_samples[25970]=26931;
squeal_samples[25971]=28991;
squeal_samples[25972]=30958;
squeal_samples[25973]=32842;
squeal_samples[25974]=34647;
squeal_samples[25975]=36354;
squeal_samples[25976]=38001;
squeal_samples[25977]=39563;
squeal_samples[25978]=41064;
squeal_samples[25979]=42490;
squeal_samples[25980]=43858;
squeal_samples[25981]=45160;
squeal_samples[25982]=46408;
squeal_samples[25983]=47598;
squeal_samples[25984]=48732;
squeal_samples[25985]=49818;
squeal_samples[25986]=50852;
squeal_samples[25987]=51839;
squeal_samples[25988]=52788;
squeal_samples[25989]=53692;
squeal_samples[25990]=53240;
squeal_samples[25991]=47951;
squeal_samples[25992]=42546;
squeal_samples[25993]=37488;
squeal_samples[25994]=32754;
squeal_samples[25995]=28315;
squeal_samples[25996]=24170;
squeal_samples[25997]=20294;
squeal_samples[25998]=16667;
squeal_samples[25999]=13261;
squeal_samples[26000]=10082;
squeal_samples[26001]=7109;
squeal_samples[26002]=5039;
squeal_samples[26003]=7363;
squeal_samples[26004]=10275;
squeal_samples[26005]=13077;
squeal_samples[26006]=15748;
squeal_samples[26007]=18301;
squeal_samples[26008]=20742;
squeal_samples[26009]=23082;
squeal_samples[26010]=25304;
squeal_samples[26011]=27444;
squeal_samples[26012]=29482;
squeal_samples[26013]=31430;
squeal_samples[26014]=33293;
squeal_samples[26015]=35065;
squeal_samples[26016]=36766;
squeal_samples[26017]=38385;
squeal_samples[26018]=39936;
squeal_samples[26019]=41413;
squeal_samples[26020]=42826;
squeal_samples[26021]=44178;
squeal_samples[26022]=45467;
squeal_samples[26023]=46697;
squeal_samples[26024]=47872;
squeal_samples[26025]=48998;
squeal_samples[26026]=50068;
squeal_samples[26027]=51094;
squeal_samples[26028]=52073;
squeal_samples[26029]=53011;
squeal_samples[26030]=53902;
squeal_samples[26031]=52183;
squeal_samples[26032]=46551;
squeal_samples[26033]=41237;
squeal_samples[26034]=36260;
squeal_samples[26035]=31606;
squeal_samples[26036]=27246;
squeal_samples[26037]=23164;
squeal_samples[26038]=19349;
squeal_samples[26039]=15780;
squeal_samples[26040]=12436;
squeal_samples[26041]=9308;
squeal_samples[26042]=6385;
squeal_samples[26043]=5258;
squeal_samples[26044]=8093;
squeal_samples[26045]=10978;
squeal_samples[26046]=13743;
squeal_samples[26047]=16383;
squeal_samples[26048]=18912;
squeal_samples[26049]=21331;
squeal_samples[26050]=23628;
squeal_samples[26051]=25843;
squeal_samples[26052]=27949;
squeal_samples[26053]=29964;
squeal_samples[26054]=31893;
squeal_samples[26055]=33727;
squeal_samples[26056]=35493;
squeal_samples[26057]=37161;
squeal_samples[26058]=38775;
squeal_samples[26059]=40299;
squeal_samples[26060]=41762;
squeal_samples[26061]=43162;
squeal_samples[26062]=44490;
squeal_samples[26063]=45766;
squeal_samples[26064]=46984;
squeal_samples[26065]=48141;
squeal_samples[26066]=49260;
squeal_samples[26067]=50315;
squeal_samples[26068]=51328;
squeal_samples[26069]=52296;
squeal_samples[26070]=53220;
squeal_samples[26071]=54059;
squeal_samples[26072]=50764;
squeal_samples[26073]=45178;
squeal_samples[26074]=39955;
squeal_samples[26075]=35051;
squeal_samples[26076]=30479;
squeal_samples[26077]=26184;
squeal_samples[26078]=22175;
squeal_samples[26079]=18420;
squeal_samples[26080]=14909;
squeal_samples[26081]=11621;
squeal_samples[26082]=8548;
squeal_samples[26083]=5669;
squeal_samples[26084]=5830;
squeal_samples[26085]=8814;
squeal_samples[26086]=11668;
squeal_samples[26087]=14399;
squeal_samples[26088]=17017;
squeal_samples[26089]=19516;
squeal_samples[26090]=21897;
squeal_samples[26091]=24185;
squeal_samples[26092]=26364;
squeal_samples[26093]=28450;
squeal_samples[26094]=30442;
squeal_samples[26095]=32345;
squeal_samples[26096]=34163;
squeal_samples[26097]=35902;
squeal_samples[26098]=37559;
squeal_samples[26099]=39147;
squeal_samples[26100]=40656;
squeal_samples[26101]=42109;
squeal_samples[26102]=43486;
squeal_samples[26103]=44804;
squeal_samples[26104]=46066;
squeal_samples[26105]=47266;
squeal_samples[26106]=48418;
squeal_samples[26107]=49514;
squeal_samples[26108]=50562;
squeal_samples[26109]=51565;
squeal_samples[26110]=52524;
squeal_samples[26111]=53439;
squeal_samples[26112]=53834;
squeal_samples[26113]=49324;
squeal_samples[26114]=43830;
squeal_samples[26115]=38687;
squeal_samples[26116]=33870;
squeal_samples[26117]=29360;
squeal_samples[26118]=25151;
squeal_samples[26119]=21203;
squeal_samples[26120]=17517;
squeal_samples[26121]=14052;
squeal_samples[26122]=10824;
squeal_samples[26123]=7795;
squeal_samples[26124]=5148;
squeal_samples[26125]=6574;
squeal_samples[26126]=9525;
squeal_samples[26127]=12351;
squeal_samples[26128]=15056;
squeal_samples[26129]=17640;
squeal_samples[26130]=20113;
squeal_samples[26131]=22466;
squeal_samples[26132]=24727;
squeal_samples[26133]=26884;
squeal_samples[26134]=28943;
squeal_samples[26135]=30917;
squeal_samples[26136]=32797;
squeal_samples[26137]=34596;
squeal_samples[26138]=36313;
squeal_samples[26139]=37948;
squeal_samples[26140]=39520;
squeal_samples[26141]=41015;
squeal_samples[26142]=42444;
squeal_samples[26143]=43811;
squeal_samples[26144]=45113;
squeal_samples[26145]=46361;
squeal_samples[26146]=47552;
squeal_samples[26147]=48683;
squeal_samples[26148]=49774;
squeal_samples[26149]=50801;
squeal_samples[26150]=51796;
squeal_samples[26151]=52739;
squeal_samples[26152]=53646;
squeal_samples[26153]=53192;
squeal_samples[26154]=47905;
squeal_samples[26155]=42498;
squeal_samples[26156]=37442;
squeal_samples[26157]=32707;
squeal_samples[26158]=28268;
squeal_samples[26159]=24122;
squeal_samples[26160]=20250;
squeal_samples[26161]=16616;
squeal_samples[26162]=13217;
squeal_samples[26163]=10036;
squeal_samples[26164]=7057;
squeal_samples[26165]=5000;
squeal_samples[26166]=7308;
squeal_samples[26167]=10233;
squeal_samples[26168]=13028;
squeal_samples[26169]=15703;
squeal_samples[26170]=18252;
squeal_samples[26171]=20698;
squeal_samples[26172]=23029;
squeal_samples[26173]=25263;
squeal_samples[26174]=27395;
squeal_samples[26175]=29435;
squeal_samples[26176]=31383;
squeal_samples[26177]=33246;
squeal_samples[26178]=35017;
squeal_samples[26179]=36720;
squeal_samples[26180]=38339;
squeal_samples[26181]=39886;
squeal_samples[26182]=41369;
squeal_samples[26183]=42777;
squeal_samples[26184]=44131;
squeal_samples[26185]=45422;
squeal_samples[26186]=46646;
squeal_samples[26187]=47829;
squeal_samples[26188]=48947;
squeal_samples[26189]=50024;
squeal_samples[26190]=51044;
squeal_samples[26191]=52029;
squeal_samples[26192]=52959;
squeal_samples[26193]=53859;
squeal_samples[26194]=52809;
squeal_samples[26195]=47297;
squeal_samples[26196]=41925;
squeal_samples[26197]=36904;
squeal_samples[26198]=32200;
squeal_samples[26199]=27801;
squeal_samples[26200]=23681;
squeal_samples[26201]=19830;
squeal_samples[26202]=16225;
squeal_samples[26203]=12851;
squeal_samples[26204]=9698;
squeal_samples[26205]=6738;
squeal_samples[26206]=5098;
squeal_samples[26207]=7719;
squeal_samples[26208]=10620;
squeal_samples[26209]=13399;
squeal_samples[26210]=16052;
squeal_samples[26211]=18596;
squeal_samples[26212]=21021;
squeal_samples[26213]=23339;
squeal_samples[26214]=25554;
squeal_samples[26215]=27676;
squeal_samples[26216]=29700;
squeal_samples[26217]=31638;
squeal_samples[26218]=33483;
squeal_samples[26219]=35251;
squeal_samples[26220]=36940;
squeal_samples[26221]=38549;
squeal_samples[26222]=40087;
squeal_samples[26223]=41558;
squeal_samples[26224]=42960;
squeal_samples[26225]=44306;
squeal_samples[26226]=45579;
squeal_samples[26227]=46808;
squeal_samples[26228]=47970;
squeal_samples[26229]=49092;
squeal_samples[26230]=50155;
squeal_samples[26231]=51170;
squeal_samples[26232]=52146;
squeal_samples[26233]=53075;
squeal_samples[26234]=53966;
squeal_samples[26235]=52234;
squeal_samples[26236]=46603;
squeal_samples[26237]=41281;
squeal_samples[26238]=36297;
squeal_samples[26239]=31638;
squeal_samples[26240]=27264;
squeal_samples[26241]=23190;
squeal_samples[26242]=19358;
squeal_samples[26243]=15793;
squeal_samples[26244]=12436;
squeal_samples[26245]=9311;
squeal_samples[26246]=6378;
squeal_samples[26247]=5249;
squeal_samples[26248]=8082;
squeal_samples[26249]=10970;
squeal_samples[26250]=13725;
squeal_samples[26251]=16371;
squeal_samples[26252]=18888;
squeal_samples[26253]=21311;
squeal_samples[26254]=23610;
squeal_samples[26255]=25817;
squeal_samples[26256]=27926;
squeal_samples[26257]=29938;
squeal_samples[26258]=31864;
squeal_samples[26259]=33706;
squeal_samples[26260]=35455;
squeal_samples[26261]=37134;
squeal_samples[26262]=38734;
squeal_samples[26263]=40264;
squeal_samples[26264]=41732;
squeal_samples[26265]=43120;
squeal_samples[26266]=44464;
squeal_samples[26267]=45724;
squeal_samples[26268]=46948;
squeal_samples[26269]=48105;
squeal_samples[26270]=49216;
squeal_samples[26271]=50272;
squeal_samples[26272]=51292;
squeal_samples[26273]=52251;
squeal_samples[26274]=53179;
squeal_samples[26275]=54062;
squeal_samples[26276]=51549;
squeal_samples[26277]=45906;
squeal_samples[26278]=40630;
squeal_samples[26279]=35681;
squeal_samples[26280]=31066;
squeal_samples[26281]=26728;
squeal_samples[26282]=22680;
squeal_samples[26283]=18896;
squeal_samples[26284]=15346;
squeal_samples[26285]=12027;
squeal_samples[26286]=8921;
squeal_samples[26287]=6015;
squeal_samples[26288]=5488;
squeal_samples[26289]=8437;
squeal_samples[26290]=11314;
squeal_samples[26291]=14049;
squeal_samples[26292]=16684;
squeal_samples[26293]=19189;
squeal_samples[26294]=21589;
squeal_samples[26295]=23882;
squeal_samples[26296]=26072;
squeal_samples[26297]=28174;
squeal_samples[26298]=30175;
squeal_samples[26299]=32088;
squeal_samples[26300]=33913;
squeal_samples[26301]=35665;
squeal_samples[26302]=37325;
squeal_samples[26303]=38919;
squeal_samples[26304]=40443;
squeal_samples[26305]=41896;
squeal_samples[26306]=43281;
squeal_samples[26307]=44610;
squeal_samples[26308]=45874;
squeal_samples[26309]=47081;
squeal_samples[26310]=48235;
squeal_samples[26311]=49339;
squeal_samples[26312]=50392;
squeal_samples[26313]=51398;
squeal_samples[26314]=52360;
squeal_samples[26315]=53283;
squeal_samples[26316]=54103;
squeal_samples[26317]=50811;
squeal_samples[26318]=45214;
squeal_samples[26319]=39981;
squeal_samples[26320]=35082;
squeal_samples[26321]=30489;
squeal_samples[26322]=26201;
squeal_samples[26323]=22176;
squeal_samples[26324]=18428;
squeal_samples[26325]=14908;
squeal_samples[26326]=11615;
squeal_samples[26327]=8538;
squeal_samples[26328]=5653;
squeal_samples[26329]=5813;
squeal_samples[26330]=8792;
squeal_samples[26331]=11647;
squeal_samples[26332]=14376;
squeal_samples[26333]=16992;
squeal_samples[26334]=19486;
squeal_samples[26335]=21866;
squeal_samples[26336]=24151;
squeal_samples[26337]=26334;
squeal_samples[26338]=28414;
squeal_samples[26339]=30407;
squeal_samples[26340]=32303;
squeal_samples[26341]=34130;
squeal_samples[26342]=35859;
squeal_samples[26343]=37519;
squeal_samples[26344]=39100;
squeal_samples[26345]=40616;
squeal_samples[26346]=42058;
squeal_samples[26347]=43439;
squeal_samples[26348]=44753;
squeal_samples[26349]=46017;
squeal_samples[26350]=47219;
squeal_samples[26351]=48366;
squeal_samples[26352]=49463;
squeal_samples[26353]=50511;
squeal_samples[26354]=51510;
squeal_samples[26355]=52471;
squeal_samples[26356]=53375;
squeal_samples[26357]=54045;
squeal_samples[26358]=50074;
squeal_samples[26359]=44536;
squeal_samples[26360]=39333;
squeal_samples[26361]=34482;
squeal_samples[26362]=29923;
squeal_samples[26363]=25673;
squeal_samples[26364]=21680;
squeal_samples[26365]=17963;
squeal_samples[26366]=14469;
squeal_samples[26367]=11211;
squeal_samples[26368]=8153;
squeal_samples[26369]=5339;
squeal_samples[26370]=6176;
squeal_samples[26371]=9145;
squeal_samples[26372]=11982;
squeal_samples[26373]=14696;
squeal_samples[26374]=17296;
squeal_samples[26375]=19778;
squeal_samples[26376]=22148;
squeal_samples[26377]=24416;
squeal_samples[26378]=26586;
squeal_samples[26379]=28656;
squeal_samples[26380]=30635;
squeal_samples[26381]=32530;
squeal_samples[26382]=34335;
squeal_samples[26383]=36064;
squeal_samples[26384]=37709;
squeal_samples[26385]=39288;
squeal_samples[26386]=40785;
squeal_samples[26387]=42229;
squeal_samples[26388]=43590;
squeal_samples[26389]=44911;
squeal_samples[26390]=46151;
squeal_samples[26391]=47359;
squeal_samples[26392]=48492;
squeal_samples[26393]=49588;
squeal_samples[26394]=50625;
squeal_samples[26395]=51617;
squeal_samples[26396]=52574;
squeal_samples[26397]=53479;
squeal_samples[26398]=53874;
squeal_samples[26399]=49353;
squeal_samples[26400]=43852;
squeal_samples[26401]=38702;
squeal_samples[26402]=33878;
squeal_samples[26403]=29369;
squeal_samples[26404]=25145;
squeal_samples[26405]=21201;
squeal_samples[26406]=17501;
squeal_samples[26407]=14043;
squeal_samples[26408]=10801;
squeal_samples[26409]=7772;
squeal_samples[26410]=5120;
squeal_samples[26411]=6546;
squeal_samples[26412]=9491;
squeal_samples[26413]=12320;
squeal_samples[26414]=15014;
squeal_samples[26415]=17604;
squeal_samples[26416]=20067;
squeal_samples[26417]=22421;
squeal_samples[26418]=24684;
squeal_samples[26419]=26833;
squeal_samples[26420]=28900;
squeal_samples[26421]=30868;
squeal_samples[26422]=32745;
squeal_samples[26423]=34542;
squeal_samples[26424]=36262;
squeal_samples[26425]=37899;
squeal_samples[26426]=39467;
squeal_samples[26427]=40956;
squeal_samples[26428]=42393;
squeal_samples[26429]=43746;
squeal_samples[26430]=45055;
squeal_samples[26431]=46294;
squeal_samples[26432]=47486;
squeal_samples[26433]=48617;
squeal_samples[26434]=49708;
squeal_samples[26435]=50741;
squeal_samples[26436]=51728;
squeal_samples[26437]=52674;
squeal_samples[26438]=53578;
squeal_samples[26439]=53594;
squeal_samples[26440]=48632;
squeal_samples[26441]=43176;
squeal_samples[26442]=38072;
squeal_samples[26443]=33291;
squeal_samples[26444]=28811;
squeal_samples[26445]=24627;
squeal_samples[26446]=20708;
squeal_samples[26447]=17047;
squeal_samples[26448]=13612;
squeal_samples[26449]=10402;
squeal_samples[26450]=7399;
squeal_samples[26451]=4992;
squeal_samples[26452]=6910;
squeal_samples[26453]=9843;
squeal_samples[26454]=12650;
squeal_samples[26455]=15335;
squeal_samples[26456]=17907;
squeal_samples[26457]=20358;
squeal_samples[26458]=22699;
squeal_samples[26459]=24947;
squeal_samples[26460]=27089;
squeal_samples[26461]=29136;
squeal_samples[26462]=31097;
squeal_samples[26463]=32960;
squeal_samples[26464]=34754;
squeal_samples[26465]=36455;
squeal_samples[26466]=38085;
squeal_samples[26467]=39641;
squeal_samples[26468]=41130;
squeal_samples[26469]=42547;
squeal_samples[26470]=43909;
squeal_samples[26471]=45196;
squeal_samples[26472]=46439;
squeal_samples[26473]=47616;
squeal_samples[26474]=48751;
squeal_samples[26475]=49822;
squeal_samples[26476]=50858;
squeal_samples[26477]=51840;
squeal_samples[26478]=52775;
squeal_samples[26479]=53679;
squeal_samples[26480]=53209;
squeal_samples[26481]=47923;
squeal_samples[26482]=42504;
squeal_samples[26483]=37448;
squeal_samples[26484]=32698;
squeal_samples[26485]=28262;
squeal_samples[26486]=24110;
squeal_samples[26487]=20224;
squeal_samples[26488]=16590;
squeal_samples[26489]=13188;
squeal_samples[26490]=10003;
squeal_samples[26491]=7025;
squeal_samples[26492]=4951;
squeal_samples[26493]=7276;
squeal_samples[26494]=10184;
squeal_samples[26495]=12979;
squeal_samples[26496]=15651;
squeal_samples[26497]=18203;
squeal_samples[26498]=20645;
squeal_samples[26499]=22977;
squeal_samples[26500]=25204;
squeal_samples[26501]=27341;
squeal_samples[26502]=29372;
squeal_samples[26503]=31323;
squeal_samples[26504]=33178;
squeal_samples[26505]=34958;
squeal_samples[26506]=36651;
squeal_samples[26507]=38272;
squeal_samples[26508]=39821;
squeal_samples[26509]=41300;
squeal_samples[26510]=42712;
squeal_samples[26511]=44058;
squeal_samples[26512]=45348;
squeal_samples[26513]=46578;
squeal_samples[26514]=47752;
squeal_samples[26515]=48874;
squeal_samples[26516]=49941;
squeal_samples[26517]=50970;
squeal_samples[26518]=51949;
squeal_samples[26519]=52877;
squeal_samples[26520]=53775;
squeal_samples[26521]=53307;
squeal_samples[26522]=48007;
squeal_samples[26523]=42587;
squeal_samples[26524]=37516;
squeal_samples[26525]=32767;
squeal_samples[26526]=28329;
squeal_samples[26527]=24164;
squeal_samples[26528]=20283;
squeal_samples[26529]=16639;
squeal_samples[26530]=13231;
squeal_samples[26531]=10044;
squeal_samples[26532]=7060;
squeal_samples[26533]=4996;
squeal_samples[26534]=7301;
squeal_samples[26535]=10219;
squeal_samples[26536]=13011;
squeal_samples[26537]=15675;
squeal_samples[26538]=18230;
squeal_samples[26539]=20673;
squeal_samples[26540]=22994;
squeal_samples[26541]=25229;
squeal_samples[26542]=27358;
squeal_samples[26543]=29395;
squeal_samples[26544]=31338;
squeal_samples[26545]=33193;
squeal_samples[26546]=34968;
squeal_samples[26547]=36667;
squeal_samples[26548]=38281;
squeal_samples[26549]=39831;
squeal_samples[26550]=41311;
squeal_samples[26551]=42721;
squeal_samples[26552]=44069;
squeal_samples[26553]=45352;
squeal_samples[26554]=46581;
squeal_samples[26555]=47758;
squeal_samples[26556]=48878;
squeal_samples[26557]=49947;
squeal_samples[26558]=50972;
squeal_samples[26559]=51951;
squeal_samples[26560]=52878;
squeal_samples[26561]=53782;
squeal_samples[26562]=53306;
squeal_samples[26563]=48004;
squeal_samples[26564]=42588;
squeal_samples[26565]=37514;
squeal_samples[26566]=32767;
squeal_samples[26567]=28327;
squeal_samples[26568]=24164;
squeal_samples[26569]=20281;
squeal_samples[26570]=16633;
squeal_samples[26571]=13232;
squeal_samples[26572]=10039;
squeal_samples[26573]=7060;
squeal_samples[26574]=4983;
squeal_samples[26575]=7300;
squeal_samples[26576]=10211;
squeal_samples[26577]=13002;
squeal_samples[26578]=15674;
squeal_samples[26579]=18219;
squeal_samples[26580]=20664;
squeal_samples[26581]=22987;
squeal_samples[26582]=25222;
squeal_samples[26583]=27346;
squeal_samples[26584]=29385;
squeal_samples[26585]=31329;
squeal_samples[26586]=33189;
squeal_samples[26587]=34960;
squeal_samples[26588]=36655;
squeal_samples[26589]=38278;
squeal_samples[26590]=39821;
squeal_samples[26591]=41301;
squeal_samples[26592]=42708;
squeal_samples[26593]=44059;
squeal_samples[26594]=45339;
squeal_samples[26595]=46577;
squeal_samples[26596]=47744;
squeal_samples[26597]=48872;
squeal_samples[26598]=49941;
squeal_samples[26599]=50962;
squeal_samples[26600]=51940;
squeal_samples[26601]=52873;
squeal_samples[26602]=53764;
squeal_samples[26603]=53299;
squeal_samples[26604]=47996;
squeal_samples[26605]=42576;
squeal_samples[26606]=37502;
squeal_samples[26607]=32758;
squeal_samples[26608]=28311;
squeal_samples[26609]=24159;
squeal_samples[26610]=20262;
squeal_samples[26611]=16628;
squeal_samples[26612]=13214;
squeal_samples[26613]=10032;
squeal_samples[26614]=7045;
squeal_samples[26615]=4974;
squeal_samples[26616]=7288;
squeal_samples[26617]=10196;
squeal_samples[26618]=12996;
squeal_samples[26619]=15655;
squeal_samples[26620]=18215;
squeal_samples[26621]=20651;
squeal_samples[26622]=22981;
squeal_samples[26623]=25206;
squeal_samples[26624]=27338;
squeal_samples[26625]=29370;
squeal_samples[26626]=31320;
squeal_samples[26627]=33176;
squeal_samples[26628]=34949;
squeal_samples[26629]=36648;
squeal_samples[26630]=38266;
squeal_samples[26631]=39811;
squeal_samples[26632]=41288;
squeal_samples[26633]=42698;
squeal_samples[26634]=44044;
squeal_samples[26635]=45336;
squeal_samples[26636]=46562;
squeal_samples[26637]=47736;
squeal_samples[26638]=48858;
squeal_samples[26639]=49931;
squeal_samples[26640]=50948;
squeal_samples[26641]=51930;
squeal_samples[26642]=52860;
squeal_samples[26643]=53754;
squeal_samples[26644]=53286;
squeal_samples[26645]=47985;
squeal_samples[26646]=42564;
squeal_samples[26647]=37491;
squeal_samples[26648]=32744;
squeal_samples[26649]=28303;
squeal_samples[26650]=24142;
squeal_samples[26651]=20256;
squeal_samples[26652]=16611;
squeal_samples[26653]=13208;
squeal_samples[26654]=10015;
squeal_samples[26655]=7037;
squeal_samples[26656]=4960;
squeal_samples[26657]=7276;
squeal_samples[26658]=10187;
squeal_samples[26659]=12981;
squeal_samples[26660]=15648;
squeal_samples[26661]=18198;
squeal_samples[26662]=20644;
squeal_samples[26663]=22965;
squeal_samples[26664]=25198;
squeal_samples[26665]=27324;
squeal_samples[26666]=29360;
squeal_samples[26667]=31308;
squeal_samples[26668]=33163;
squeal_samples[26669]=34940;
squeal_samples[26670]=36634;
squeal_samples[26671]=38256;
squeal_samples[26672]=39798;
squeal_samples[26673]=41277;
squeal_samples[26674]=42686;
squeal_samples[26675]=44033;
squeal_samples[26676]=45323;
squeal_samples[26677]=46554;
squeal_samples[26678]=47719;
squeal_samples[26679]=48851;
squeal_samples[26680]=49915;
squeal_samples[26681]=50940;
squeal_samples[26682]=51918;
squeal_samples[26683]=52847;
squeal_samples[26684]=53744;
squeal_samples[26685]=53272;
squeal_samples[26686]=47976;
squeal_samples[26687]=42550;
squeal_samples[26688]=37481;
squeal_samples[26689]=32731;
squeal_samples[26690]=28294;
squeal_samples[26691]=24127;
squeal_samples[26692]=20248;
squeal_samples[26693]=16595;
squeal_samples[26694]=13199;
squeal_samples[26695]=10004;
squeal_samples[26696]=7024;
squeal_samples[26697]=4950;
squeal_samples[26698]=7262;
squeal_samples[26699]=10178;
squeal_samples[26700]=12967;
squeal_samples[26701]=15638;
squeal_samples[26702]=18186;
squeal_samples[26703]=20632;
squeal_samples[26704]=22954;
squeal_samples[26705]=25185;
squeal_samples[26706]=27314;
squeal_samples[26707]=29347;
squeal_samples[26708]=31297;
squeal_samples[26709]=33151;
squeal_samples[26710]=34928;
squeal_samples[26711]=36624;
squeal_samples[26712]=38242;
squeal_samples[26713]=39789;
squeal_samples[26714]=41263;
squeal_samples[26715]=42676;
squeal_samples[26716]=44020;
squeal_samples[26717]=45314;
squeal_samples[26718]=46538;
squeal_samples[26719]=47712;
squeal_samples[26720]=48836;
squeal_samples[26721]=49905;
squeal_samples[26722]=50929;
squeal_samples[26723]=51905;
squeal_samples[26724]=52836;
squeal_samples[26725]=53731;
squeal_samples[26726]=53262;
squeal_samples[26727]=47964;
squeal_samples[26728]=42539;
squeal_samples[26729]=37469;
squeal_samples[26730]=32719;
squeal_samples[26731]=28281;
squeal_samples[26732]=24119;
squeal_samples[26733]=20232;
squeal_samples[26734]=16589;
squeal_samples[26735]=13181;
squeal_samples[26736]=9998;
squeal_samples[26737]=7008;
squeal_samples[26738]=4941;
squeal_samples[26739]=7250;
squeal_samples[26740]=10165;
squeal_samples[26741]=12958;
squeal_samples[26742]=15624;
squeal_samples[26743]=18176;
squeal_samples[26744]=20619;
squeal_samples[26745]=22944;
squeal_samples[26746]=25172;
squeal_samples[26747]=27304;
squeal_samples[26748]=29334;
squeal_samples[26749]=31287;
squeal_samples[26750]=33138;
squeal_samples[26751]=34917;
squeal_samples[26752]=36612;
squeal_samples[26753]=38232;
squeal_samples[26754]=39774;
squeal_samples[26755]=41256;
squeal_samples[26756]=42660;
squeal_samples[26757]=44012;
squeal_samples[26758]=45300;
squeal_samples[26759]=46526;
squeal_samples[26760]=47703;
squeal_samples[26761]=48822;
squeal_samples[26762]=49896;
squeal_samples[26763]=50913;
squeal_samples[26764]=51896;
squeal_samples[26765]=52825;
squeal_samples[26766]=53718;
squeal_samples[26767]=53253;
squeal_samples[26768]=47948;
squeal_samples[26769]=42530;
squeal_samples[26770]=37457;
squeal_samples[26771]=32708;
squeal_samples[26772]=28268;
squeal_samples[26773]=24109;
squeal_samples[26774]=20219;
squeal_samples[26775]=16577;
squeal_samples[26776]=13172;
squeal_samples[26777]=9982;
squeal_samples[26778]=7000;
squeal_samples[26779]=4928;
squeal_samples[26780]=7238;
squeal_samples[26781]=10155;
squeal_samples[26782]=12943;
squeal_samples[26783]=15615;
squeal_samples[26784]=18163;
squeal_samples[26785]=20609;
squeal_samples[26786]=22931;
squeal_samples[26787]=25161;
squeal_samples[26788]=27291;
squeal_samples[26789]=29324;
squeal_samples[26790]=31274;
squeal_samples[26791]=33128;
squeal_samples[26792]=34904;
squeal_samples[26793]=36601;
squeal_samples[26794]=38219;
squeal_samples[26795]=39766;
squeal_samples[26796]=41239;
squeal_samples[26797]=42654;
squeal_samples[26798]=43995;
squeal_samples[26799]=45293;
squeal_samples[26800]=46512;
squeal_samples[26801]=47692;
squeal_samples[26802]=48809;
squeal_samples[26803]=49885;
squeal_samples[26804]=50903;
squeal_samples[26805]=51883;
squeal_samples[26806]=52814;
squeal_samples[26807]=53706;
squeal_samples[26808]=53240;
squeal_samples[26809]=47939;
squeal_samples[26810]=42517;
squeal_samples[26811]=37446;
squeal_samples[26812]=32696;
squeal_samples[26813]=28256;
squeal_samples[26814]=24098;
squeal_samples[26815]=20206;
squeal_samples[26816]=16569;
squeal_samples[26817]=13156;
squeal_samples[26818]=9974;
squeal_samples[26819]=6986;
squeal_samples[26820]=4917;
squeal_samples[26821]=7227;
squeal_samples[26822]=10143;
squeal_samples[26823]=12933;
squeal_samples[26824]=15601;
squeal_samples[26825]=18153;
squeal_samples[26826]=20596;
squeal_samples[26827]=22920;
squeal_samples[26828]=25151;
squeal_samples[26829]=27277;
squeal_samples[26830]=29314;
squeal_samples[26831]=31260;
squeal_samples[26832]=33118;
squeal_samples[26833]=34893;
squeal_samples[26834]=36587;
squeal_samples[26835]=38210;
squeal_samples[26836]=39751;
squeal_samples[26837]=41230;
squeal_samples[26838]=42641;
squeal_samples[26839]=43984;
squeal_samples[26840]=45280;
squeal_samples[26841]=46502;
squeal_samples[26842]=47679;
squeal_samples[26843]=48799;
squeal_samples[26844]=49871;
squeal_samples[26845]=50894;
squeal_samples[26846]=51867;
squeal_samples[26847]=52805;
squeal_samples[26848]=53692;
squeal_samples[26849]=53702;
squeal_samples[26850]=48725;
squeal_samples[26851]=43255;
squeal_samples[26852]=38139;
squeal_samples[26853]=33343;
squeal_samples[26854]=28858;
squeal_samples[26855]=24660;
squeal_samples[26856]=20734;
squeal_samples[26857]=17060;
squeal_samples[26858]=13613;
squeal_samples[26859]=10403;
squeal_samples[26860]=7385;
squeal_samples[26861]=4979;
squeal_samples[26862]=6886;
squeal_samples[26863]=9823;
squeal_samples[26864]=12615;
squeal_samples[26865]=15305;
squeal_samples[26866]=17860;
squeal_samples[26867]=20323;
squeal_samples[26868]=22655;
squeal_samples[26869]=24901;
squeal_samples[26870]=27038;
squeal_samples[26871]=29084;
squeal_samples[26872]=31039;
squeal_samples[26873]=32904;
squeal_samples[26874]=34692;
squeal_samples[26875]=36390;
squeal_samples[26876]=38026;
squeal_samples[26877]=39569;
squeal_samples[26878]=41065;
squeal_samples[26879]=42472;
squeal_samples[26880]=43837;
squeal_samples[26881]=45122;
squeal_samples[26882]=46365;
squeal_samples[26883]=47538;
squeal_samples[26884]=48666;
squeal_samples[26885]=49737;
squeal_samples[26886]=50775;
squeal_samples[26887]=51748;
squeal_samples[26888]=52693;
squeal_samples[26889]=53589;
squeal_samples[26890]=53972;
squeal_samples[26891]=49436;
squeal_samples[26892]=43918;
squeal_samples[26893]=38757;
squeal_samples[26894]=33923;
squeal_samples[26895]=29400;
squeal_samples[26896]=25166;
squeal_samples[26897]=21203;
squeal_samples[26898]=17507;
squeal_samples[26899]=14028;
squeal_samples[26900]=10789;
squeal_samples[26901]=7744;
squeal_samples[26902]=5090;
squeal_samples[26903]=6508;
squeal_samples[26904]=9449;
squeal_samples[26905]=12270;
squeal_samples[26906]=14964;
squeal_samples[26907]=17544;
squeal_samples[26908]=20012;
squeal_samples[26909]=22367;
squeal_samples[26910]=24613;
squeal_samples[26911]=26770;
squeal_samples[26912]=28822;
squeal_samples[26913]=30792;
squeal_samples[26914]=32674;
squeal_samples[26915]=34456;
squeal_samples[26916]=36181;
squeal_samples[26917]=37812;
squeal_samples[26918]=39378;
squeal_samples[26919]=40870;
squeal_samples[26920]=42296;
squeal_samples[26921]=43659;
squeal_samples[26922]=44956;
squeal_samples[26923]=46199;
squeal_samples[26924]=47386;
squeal_samples[26925]=48519;
squeal_samples[26926]=49601;
squeal_samples[26927]=50637;
squeal_samples[26928]=51623;
squeal_samples[26929]=52566;
squeal_samples[26930]=53470;
squeal_samples[26931]=54122;
squeal_samples[26932]=50142;
squeal_samples[26933]=44581;
squeal_samples[26934]=39373;
squeal_samples[26935]=34501;
squeal_samples[26936]=29935;
squeal_samples[26937]=25669;
squeal_samples[26938]=21674;
squeal_samples[26939]=17940;
squeal_samples[26940]=14441;
squeal_samples[26941]=11168;
squeal_samples[26942]=8106;
squeal_samples[26943]=5283;
squeal_samples[26944]=6117;
squeal_samples[26945]=9077;
squeal_samples[26946]=11919;
squeal_samples[26947]=14622;
squeal_samples[26948]=17221;
squeal_samples[26949]=19695;
squeal_samples[26950]=22067;
squeal_samples[26951]=24328;
squeal_samples[26952]=26494;
squeal_samples[26953]=28562;
squeal_samples[26954]=30537;
squeal_samples[26955]=32427;
squeal_samples[26956]=34231;
squeal_samples[26957]=35955;
squeal_samples[26958]=37600;
squeal_samples[26959]=39173;
squeal_samples[26960]=40671;
squeal_samples[26961]=42109;
squeal_samples[26962]=43476;
squeal_samples[26963]=44790;
squeal_samples[26964]=46032;
squeal_samples[26965]=47231;
squeal_samples[26966]=48370;
squeal_samples[26967]=49455;
squeal_samples[26968]=50499;
squeal_samples[26969]=51487;
squeal_samples[26970]=52440;
squeal_samples[26971]=53344;
squeal_samples[26972]=54164;
squeal_samples[26973]=50848;
squeal_samples[26974]=45243;
squeal_samples[26975]=39992;
squeal_samples[26976]=35081;
squeal_samples[26977]=30476;
squeal_samples[26978]=26182;
squeal_samples[26979]=22147;
squeal_samples[26980]=18382;
squeal_samples[26981]=14857;
squeal_samples[26982]=11554;
squeal_samples[26983]=8469;
squeal_samples[26984]=5577;
squeal_samples[26985]=5727;
squeal_samples[26986]=8706;
squeal_samples[26987]=11555;
squeal_samples[26988]=14284;
squeal_samples[26989]=16890;
squeal_samples[26990]=19383;
squeal_samples[26991]=21760;
squeal_samples[26992]=24041;
squeal_samples[26993]=26215;
squeal_samples[26994]=28296;
squeal_samples[26995]=30288;
squeal_samples[26996]=32185;
squeal_samples[26997]=34001;
squeal_samples[26998]=35726;
squeal_samples[26999]=37394;
squeal_samples[27000]=38965;
squeal_samples[27001]=40482;
squeal_samples[27002]=41917;
squeal_samples[27003]=43302;
squeal_samples[27004]=44611;
squeal_samples[27005]=45872;
squeal_samples[27006]=47072;
squeal_samples[27007]=48215;
squeal_samples[27008]=49317;
squeal_samples[27009]=50352;
squeal_samples[27010]=51361;
squeal_samples[27011]=52306;
squeal_samples[27012]=53224;
squeal_samples[27013]=54097;
squeal_samples[27014]=51567;
squeal_samples[27015]=45912;
squeal_samples[27016]=40621;
squeal_samples[27017]=35661;
squeal_samples[27018]=31030;
squeal_samples[27019]=26687;
squeal_samples[27020]=22627;
squeal_samples[27021]=18830;
squeal_samples[27022]=15271;
squeal_samples[27023]=11942;
squeal_samples[27024]=8836;
squeal_samples[27025]=5915;
squeal_samples[27026]=5381;
squeal_samples[27027]=8329;
squeal_samples[27028]=11190;
squeal_samples[27029]=13937;
squeal_samples[27030]=16557;
squeal_samples[27031]=19067;
squeal_samples[27032]=21457;
squeal_samples[27033]=23744;
squeal_samples[27034]=25942;
squeal_samples[27035]=28027;
squeal_samples[27036]=30032;
squeal_samples[27037]=31942;
squeal_samples[27038]=33763;
squeal_samples[27039]=35507;
squeal_samples[27040]=37175;
squeal_samples[27041]=38759;
squeal_samples[27042]=40284;
squeal_samples[27043]=41733;
squeal_samples[27044]=43122;
squeal_samples[27045]=44441;
squeal_samples[27046]=45711;
squeal_samples[27047]=46911;
squeal_samples[27048]=48065;
squeal_samples[27049]=49167;
squeal_samples[27050]=50218;
squeal_samples[27051]=51222;
squeal_samples[27052]=52182;
squeal_samples[27053]=53098;
squeal_samples[27054]=53976;
squeal_samples[27055]=52233;
squeal_samples[27056]=46588;
squeal_samples[27057]=41253;
squeal_samples[27058]=36255;
squeal_samples[27059]=31583;
squeal_samples[27060]=27199;
squeal_samples[27061]=23107;
squeal_samples[27062]=19280;
squeal_samples[27063]=15692;
squeal_samples[27064]=12336;
squeal_samples[27065]=9194;
squeal_samples[27066]=6262;
squeal_samples[27067]=5122;
squeal_samples[27068]=7955;
squeal_samples[27069]=10829;
squeal_samples[27070]=13590;
squeal_samples[27071]=16225;
squeal_samples[27072]=18746;
squeal_samples[27073]=21158;
squeal_samples[27074]=23455;
squeal_samples[27075]=25660;
squeal_samples[27076]=27759;
squeal_samples[27077]=29777;
squeal_samples[27078]=31697;
squeal_samples[27079]=33530;
squeal_samples[27080]=35283;
squeal_samples[27081]=36962;
squeal_samples[27082]=38553;
squeal_samples[27083]=40088;
squeal_samples[27084]=41542;
squeal_samples[27085]=42943;
squeal_samples[27086]=44267;
squeal_samples[27087]=45541;
squeal_samples[27088]=46754;
squeal_samples[27089]=47912;
squeal_samples[27090]=49018;
squeal_samples[27091]=50080;
squeal_samples[27092]=51088;
squeal_samples[27093]=52052;
squeal_samples[27094]=52977;
squeal_samples[27095]=53860;
squeal_samples[27096]=52799;
squeal_samples[27097]=47266;
squeal_samples[27098]=41888;
squeal_samples[27099]=36853;
squeal_samples[27100]=32131;
squeal_samples[27101]=27728;
squeal_samples[27102]=23587;
squeal_samples[27103]=19736;
squeal_samples[27104]=16111;
squeal_samples[27105]=12733;
squeal_samples[27106]=9564;
squeal_samples[27107]=6601;
squeal_samples[27108]=4957;
squeal_samples[27109]=7568;
squeal_samples[27110]=10471;
squeal_samples[27111]=13235;
squeal_samples[27112]=15892;
squeal_samples[27113]=18423;
squeal_samples[27114]=20853;
squeal_samples[27115]=23165;
squeal_samples[27116]=25377;
squeal_samples[27117]=27497;
squeal_samples[27118]=29513;
squeal_samples[27119]=31448;
squeal_samples[27120]=33291;
squeal_samples[27121]=35055;
squeal_samples[27122]=36742;
squeal_samples[27123]=38349;
squeal_samples[27124]=39883;
squeal_samples[27125]=41357;
squeal_samples[27126]=42752;
squeal_samples[27127]=44096;
squeal_samples[27128]=45371;
squeal_samples[27129]=46590;
squeal_samples[27130]=47760;
squeal_samples[27131]=48872;
squeal_samples[27132]=49934;
squeal_samples[27133]=50955;
squeal_samples[27134]=51925;
squeal_samples[27135]=52850;
squeal_samples[27136]=53742;
squeal_samples[27137]=53264;
squeal_samples[27138]=47955;
squeal_samples[27139]=42529;
squeal_samples[27140]=37449;
squeal_samples[27141]=32696;
squeal_samples[27142]=28247;
squeal_samples[27143]=24079;
squeal_samples[27144]=20192;
squeal_samples[27145]=16544;
squeal_samples[27146]=13130;
squeal_samples[27147]=9941;
squeal_samples[27148]=6948;
squeal_samples[27149]=4879;
squeal_samples[27150]=7183;
squeal_samples[27151]=10098;
squeal_samples[27152]=12885;
squeal_samples[27153]=15552;
squeal_samples[27154]=18103;
squeal_samples[27155]=20543;
squeal_samples[27156]=22863;
squeal_samples[27157]=25099;
squeal_samples[27158]=27220;
squeal_samples[27159]=29262;
squeal_samples[27160]=31198;
squeal_samples[27161]=33060;
squeal_samples[27162]=34830;
squeal_samples[27163]=36526;
squeal_samples[27164]=38141;
squeal_samples[27165]=39687;
squeal_samples[27166]=41166;
squeal_samples[27167]=42566;
squeal_samples[27168]=43924;
squeal_samples[27169]=45198;
squeal_samples[27170]=46437;
squeal_samples[27171]=47602;
squeal_samples[27172]=48728;
squeal_samples[27173]=49791;
squeal_samples[27174]=50818;
squeal_samples[27175]=51793;
squeal_samples[27176]=52725;
squeal_samples[27177]=53619;
squeal_samples[27178]=53991;
squeal_samples[27179]=49456;
squeal_samples[27180]=43933;
squeal_samples[27181]=38763;
squeal_samples[27182]=33924;
squeal_samples[27183]=29395;
squeal_samples[27184]=25155;
squeal_samples[27185]=21190;
squeal_samples[27186]=17482;
squeal_samples[27187]=14005;
squeal_samples[27188]=10760;
squeal_samples[27189]=7718;
squeal_samples[27190]=5059;
squeal_samples[27191]=6468;
squeal_samples[27192]=9414;
squeal_samples[27193]=12233;
squeal_samples[27194]=14924;
squeal_samples[27195]=17503;
squeal_samples[27196]=19962;
squeal_samples[27197]=22319;
squeal_samples[27198]=24567;
squeal_samples[27199]=26719;
squeal_samples[27200]=28775;
squeal_samples[27201]=30738;
squeal_samples[27202]=32619;
squeal_samples[27203]=34406;
squeal_samples[27204]=36123;
squeal_samples[27205]=37756;
squeal_samples[27206]=39317;
squeal_samples[27207]=40812;
squeal_samples[27208]=42231;
squeal_samples[27209]=43595;
squeal_samples[27210]=44896;
squeal_samples[27211]=46134;
squeal_samples[27212]=47323;
squeal_samples[27213]=48453;
squeal_samples[27214]=49537;
squeal_samples[27215]=50571;
squeal_samples[27216]=51555;
squeal_samples[27217]=52499;
squeal_samples[27218]=53401;
squeal_samples[27219]=54207;
squeal_samples[27220]=50894;
squeal_samples[27221]=45277;
squeal_samples[27222]=40020;
squeal_samples[27223]=35104;
squeal_samples[27224]=30494;
squeal_samples[27225]=26188;
squeal_samples[27226]=22149;
squeal_samples[27227]=18384;
squeal_samples[27228]=14852;
squeal_samples[27229]=11545;
squeal_samples[27230]=8453;
squeal_samples[27231]=5563;
squeal_samples[27232]=5706;
squeal_samples[27233]=8687;
squeal_samples[27234]=11526;
squeal_samples[27235]=14262;
squeal_samples[27236]=16862;
squeal_samples[27237]=19352;
squeal_samples[27238]=21728;
squeal_samples[27239]=24011;
squeal_samples[27240]=26183;
squeal_samples[27241]=28266;
squeal_samples[27242]=30249;
squeal_samples[27243]=32145;
squeal_samples[27244]=33962;
squeal_samples[27245]=35693;
squeal_samples[27246]=37348;
squeal_samples[27247]=38926;
squeal_samples[27248]=40437;
squeal_samples[27249]=41872;
squeal_samples[27250]=43253;
squeal_samples[27251]=44564;
squeal_samples[27252]=45824;
squeal_samples[27253]=47024;
squeal_samples[27254]=48169;
squeal_samples[27255]=49261;
squeal_samples[27256]=50303;
squeal_samples[27257]=51304;
squeal_samples[27258]=52254;
squeal_samples[27259]=53171;
squeal_samples[27260]=54043;
squeal_samples[27261]=52290;
squeal_samples[27262]=46639;
squeal_samples[27263]=41292;
squeal_samples[27264]=36290;
squeal_samples[27265]=31611;
squeal_samples[27266]=27225;
squeal_samples[27267]=23130;
squeal_samples[27268]=19292;
squeal_samples[27269]=15701;
squeal_samples[27270]=12341;
squeal_samples[27271]=9199;
squeal_samples[27272]=6255;
squeal_samples[27273]=5117;
squeal_samples[27274]=7942;
squeal_samples[27275]=10818;
squeal_samples[27276]=13579;
squeal_samples[27277]=16212;
squeal_samples[27278]=18731;
squeal_samples[27279]=21138;
squeal_samples[27280]=23437;
squeal_samples[27281]=25636;
squeal_samples[27282]=27745;
squeal_samples[27283]=29748;
squeal_samples[27284]=31674;
squeal_samples[27285]=33498;
squeal_samples[27286]=35253;
squeal_samples[27287]=36930;
squeal_samples[27288]=38525;
squeal_samples[27289]=40055;
squeal_samples[27290]=41509;
squeal_samples[27291]=42903;
squeal_samples[27292]=44234;
squeal_samples[27293]=45503;
squeal_samples[27294]=46714;
squeal_samples[27295]=47875;
squeal_samples[27296]=48978;
squeal_samples[27297]=50037;
squeal_samples[27298]=51046;
squeal_samples[27299]=52013;
squeal_samples[27300]=52932;
squeal_samples[27301]=53816;
squeal_samples[27302]=53331;
squeal_samples[27303]=48018;
squeal_samples[27304]=42586;
squeal_samples[27305]=37500;
squeal_samples[27306]=32740;
squeal_samples[27307]=28282;
squeal_samples[27308]=24119;
squeal_samples[27309]=20212;
squeal_samples[27310]=16572;
squeal_samples[27311]=13142;
squeal_samples[27312]=9956;
squeal_samples[27313]=6960;
squeal_samples[27314]=4888;
squeal_samples[27315]=7191;
squeal_samples[27316]=10101;
squeal_samples[27317]=12888;
squeal_samples[27318]=15549;
squeal_samples[27319]=18101;
squeal_samples[27320]=20535;
squeal_samples[27321]=22855;
squeal_samples[27322]=25084;
squeal_samples[27323]=27209;
squeal_samples[27324]=29245;
squeal_samples[27325]=31190;
squeal_samples[27326]=33036;
squeal_samples[27327]=34815;
squeal_samples[27328]=36504;
squeal_samples[27329]=38123;
squeal_samples[27330]=39665;
squeal_samples[27331]=41137;
squeal_samples[27332]=42554;
squeal_samples[27333]=43893;
squeal_samples[27334]=45179;
squeal_samples[27335]=46403;
squeal_samples[27336]=47576;
squeal_samples[27337]=48695;
squeal_samples[27338]=49764;
squeal_samples[27339]=50787;
squeal_samples[27340]=51763;
squeal_samples[27341]=52697;
squeal_samples[27342]=53587;
squeal_samples[27343]=53963;
squeal_samples[27344]=49420;
squeal_samples[27345]=43898;
squeal_samples[27346]=38728;
squeal_samples[27347]=33889;
squeal_samples[27348]=29360;
squeal_samples[27349]=25119;
squeal_samples[27350]=21151;
squeal_samples[27351]=17445;
squeal_samples[27352]=13973;
squeal_samples[27353]=10715;
squeal_samples[27354]=7683;
squeal_samples[27355]=5013;
squeal_samples[27356]=6433;
squeal_samples[27357]=9370;
squeal_samples[27358]=12193;
squeal_samples[27359]=14884;
squeal_samples[27360]=17462;
squeal_samples[27361]=19923;
squeal_samples[27362]=22278;
squeal_samples[27363]=24526;
squeal_samples[27364]=26678;
squeal_samples[27365]=28735;
squeal_samples[27366]=30697;
squeal_samples[27367]=32575;
squeal_samples[27368]=34363;
squeal_samples[27369]=36079;
squeal_samples[27370]=37715;
squeal_samples[27371]=39270;
squeal_samples[27372]=40767;
squeal_samples[27373]=42190;
squeal_samples[27374]=43555;
squeal_samples[27375]=44850;
squeal_samples[27376]=46094;
squeal_samples[27377]=47276;
squeal_samples[27378]=48412;
squeal_samples[27379]=49492;
squeal_samples[27380]=50526;
squeal_samples[27381]=51511;
squeal_samples[27382]=52458;
squeal_samples[27383]=53350;
squeal_samples[27384]=54170;
squeal_samples[27385]=50848;
squeal_samples[27386]=45234;
squeal_samples[27387]=39977;
squeal_samples[27388]=35056;
squeal_samples[27389]=30450;
squeal_samples[27390]=26140;
squeal_samples[27391]=22111;
squeal_samples[27392]=18336;
squeal_samples[27393]=14808;
squeal_samples[27394]=11497;
squeal_samples[27395]=8410;
squeal_samples[27396]=5513;
squeal_samples[27397]=5666;
squeal_samples[27398]=8634;
squeal_samples[27399]=11488;
squeal_samples[27400]=14209;
squeal_samples[27401]=16821;
squeal_samples[27402]=19309;
squeal_samples[27403]=21684;
squeal_samples[27404]=23963;
squeal_samples[27405]=26140;
squeal_samples[27406]=28218;
squeal_samples[27407]=30204;
squeal_samples[27408]=32099;
squeal_samples[27409]=33915;
squeal_samples[27410]=35649;
squeal_samples[27411]=37301;
squeal_samples[27412]=38881;
squeal_samples[27413]=40389;
squeal_samples[27414]=41829;
squeal_samples[27415]=43205;
squeal_samples[27416]=44519;
squeal_samples[27417]=45778;
squeal_samples[27418]=46977;
squeal_samples[27419]=48126;
squeal_samples[27420]=49212;
squeal_samples[27421]=50260;
squeal_samples[27422]=51256;
squeal_samples[27423]=52210;
squeal_samples[27424]=53125;
squeal_samples[27425]=53995;
squeal_samples[27426]=52248;
squeal_samples[27427]=46588;
squeal_samples[27428]=41251;
squeal_samples[27429]=36241;
squeal_samples[27430]=31566;
squeal_samples[27431]=27181;
squeal_samples[27432]=23080;
squeal_samples[27433]=19250;
squeal_samples[27434]=15651;
squeal_samples[27435]=12301;
squeal_samples[27436]=9147;
squeal_samples[27437]=6216;
squeal_samples[27438]=5064;
squeal_samples[27439]=7902;
squeal_samples[27440]=10770;
squeal_samples[27441]=13534;
squeal_samples[27442]=16165;
squeal_samples[27443]=18687;
squeal_samples[27444]=21096;
squeal_samples[27445]=23392;
squeal_samples[27446]=25592;
squeal_samples[27447]=27696;
squeal_samples[27448]=29704;
squeal_samples[27449]=31628;
squeal_samples[27450]=33451;
squeal_samples[27451]=35210;
squeal_samples[27452]=36881;
squeal_samples[27453]=38481;
squeal_samples[27454]=40009;
squeal_samples[27455]=41463;
squeal_samples[27456]=42857;
squeal_samples[27457]=44189;
squeal_samples[27458]=45456;
squeal_samples[27459]=46669;
squeal_samples[27460]=47830;
squeal_samples[27461]=48929;
squeal_samples[27462]=49994;
squeal_samples[27463]=51000;
squeal_samples[27464]=51964;
squeal_samples[27465]=52891;
squeal_samples[27466]=53765;
squeal_samples[27467]=53288;
squeal_samples[27468]=47973;
squeal_samples[27469]=42538;
squeal_samples[27470]=37455;
squeal_samples[27471]=32694;
squeal_samples[27472]=28237;
squeal_samples[27473]=24072;
squeal_samples[27474]=20169;
squeal_samples[27475]=16522;
squeal_samples[27476]=13101;
squeal_samples[27477]=9905;
squeal_samples[27478]=6918;
squeal_samples[27479]=4839;
squeal_samples[27480]=7148;
squeal_samples[27481]=10053;
squeal_samples[27482]=12844;
squeal_samples[27483]=15501;
squeal_samples[27484]=18056;
squeal_samples[27485]=20490;
squeal_samples[27486]=22807;
squeal_samples[27487]=25041;
squeal_samples[27488]=27161;
squeal_samples[27489]=29200;
squeal_samples[27490]=31144;
squeal_samples[27491]=32990;
squeal_samples[27492]=34769;
squeal_samples[27493]=36458;
squeal_samples[27494]=38078;
squeal_samples[27495]=39617;
squeal_samples[27496]=41094;
squeal_samples[27497]=42504;
squeal_samples[27498]=43850;
squeal_samples[27499]=45132;
squeal_samples[27500]=46356;
squeal_samples[27501]=47533;
squeal_samples[27502]=48645;
squeal_samples[27503]=49721;
squeal_samples[27504]=50738;
squeal_samples[27505]=51720;
squeal_samples[27506]=52648;
squeal_samples[27507]=53542;
squeal_samples[27508]=54183;
squeal_samples[27509]=50187;
squeal_samples[27510]=44615;
squeal_samples[27511]=39392;
squeal_samples[27512]=34512;
squeal_samples[27513]=29938;
squeal_samples[27514]=25659;
squeal_samples[27515]=21653;
squeal_samples[27516]=17910;
squeal_samples[27517]=14405;
squeal_samples[27518]=11120;
squeal_samples[27519]=8054;
squeal_samples[27520]=5225;
squeal_samples[27521]=6053;
squeal_samples[27522]=9009;
squeal_samples[27523]=11843;
squeal_samples[27524]=14545;
squeal_samples[27525]=17139;
squeal_samples[27526]=19612;
squeal_samples[27527]=21975;
squeal_samples[27528]=24237;
squeal_samples[27529]=26399;
squeal_samples[27530]=28466;
squeal_samples[27531]=30440;
squeal_samples[27532]=32327;
squeal_samples[27533]=34124;
squeal_samples[27534]=35846;
squeal_samples[27535]=37491;
squeal_samples[27536]=39056;
squeal_samples[27537]=40565;
squeal_samples[27538]=41990;
squeal_samples[27539]=43364;
squeal_samples[27540]=44661;
squeal_samples[27541]=45914;
squeal_samples[27542]=47105;
squeal_samples[27543]=48241;
squeal_samples[27544]=49327;
squeal_samples[27545]=50369;
squeal_samples[27546]=51360;
squeal_samples[27547]=52303;
squeal_samples[27548]=53217;
squeal_samples[27549]=54075;
squeal_samples[27550]=52325;
squeal_samples[27551]=46661;
squeal_samples[27552]=41309;
squeal_samples[27553]=36304;
squeal_samples[27554]=31613;
squeal_samples[27555]=27232;
squeal_samples[27556]=23120;
squeal_samples[27557]=19287;
squeal_samples[27558]=15688;
squeal_samples[27559]=12322;
squeal_samples[27560]=9177;
squeal_samples[27561]=6232;
squeal_samples[27562]=5087;
squeal_samples[27563]=7915;
squeal_samples[27564]=10783;
squeal_samples[27565]=13545;
squeal_samples[27566]=16173;
squeal_samples[27567]=18691;
squeal_samples[27568]=21093;
squeal_samples[27569]=23397;
squeal_samples[27570]=25594;
squeal_samples[27571]=27694;
squeal_samples[27572]=29705;
squeal_samples[27573]=31616;
squeal_samples[27574]=33455;
squeal_samples[27575]=35203;
squeal_samples[27576]=36877;
squeal_samples[27577]=38471;
squeal_samples[27578]=39998;
squeal_samples[27579]=41454;
squeal_samples[27580]=42847;
squeal_samples[27581]=44173;
squeal_samples[27582]=45446;
squeal_samples[27583]=46653;
squeal_samples[27584]=47813;
squeal_samples[27585]=48917;
squeal_samples[27586]=49975;
squeal_samples[27587]=50981;
squeal_samples[27588]=51946;
squeal_samples[27589]=52867;
squeal_samples[27590]=53746;
squeal_samples[27591]=53744;
squeal_samples[27592]=48750;
squeal_samples[27593]=43267;
squeal_samples[27594]=38131;
squeal_samples[27595]=33327;
squeal_samples[27596]=28828;
squeal_samples[27597]=24618;
squeal_samples[27598]=20682;
squeal_samples[27599]=17000;
squeal_samples[27600]=13547;
squeal_samples[27601]=10319;
squeal_samples[27602]=7301;
squeal_samples[27603]=4881;
squeal_samples[27604]=6786;
squeal_samples[27605]=9710;
squeal_samples[27606]=12509;
squeal_samples[27607]=15187;
squeal_samples[27608]=17748;
squeal_samples[27609]=20201;
squeal_samples[27610]=22528;
squeal_samples[27611]=24773;
squeal_samples[27612]=26905;
squeal_samples[27613]=28948;
squeal_samples[27614]=30903;
squeal_samples[27615]=32760;
squeal_samples[27616]=34545;
squeal_samples[27617]=36245;
squeal_samples[27618]=37870;
squeal_samples[27619]=39418;
squeal_samples[27620]=40905;
squeal_samples[27621]=42316;
squeal_samples[27622]=43671;
squeal_samples[27623]=44960;
squeal_samples[27624]=46193;
squeal_samples[27625]=47371;
squeal_samples[27626]=48501;
squeal_samples[27627]=49569;
squeal_samples[27628]=50598;
squeal_samples[27629]=51580;
squeal_samples[27630]=52515;
squeal_samples[27631]=53412;
squeal_samples[27632]=54210;
squeal_samples[27633]=50896;
squeal_samples[27634]=45267;
squeal_samples[27635]=40007;
squeal_samples[27636]=35078;
squeal_samples[27637]=30470;
squeal_samples[27638]=26150;
squeal_samples[27639]=22114;
squeal_samples[27640]=18339;
squeal_samples[27641]=14801;
squeal_samples[27642]=11498;
squeal_samples[27643]=8395;
squeal_samples[27644]=5505;
squeal_samples[27645]=5646;
squeal_samples[27646]=8619;
squeal_samples[27647]=11463;
squeal_samples[27648]=14188;
squeal_samples[27649]=16792;
squeal_samples[27650]=19283;
squeal_samples[27651]=21654;
squeal_samples[27652]=23936;
squeal_samples[27653]=26099;
squeal_samples[27654]=28187;
squeal_samples[27655]=30165;
squeal_samples[27656]=32064;
squeal_samples[27657]=33873;
squeal_samples[27658]=35607;
squeal_samples[27659]=37259;
squeal_samples[27660]=38842;
squeal_samples[27661]=40339;
squeal_samples[27662]=41789;
squeal_samples[27663]=43157;
squeal_samples[27664]=44472;
squeal_samples[27665]=45727;
squeal_samples[27666]=46923;
squeal_samples[27667]=48073;
squeal_samples[27668]=49160;
squeal_samples[27669]=50208;
squeal_samples[27670]=51202;
squeal_samples[27671]=52159;
squeal_samples[27672]=53069;
squeal_samples[27673]=53940;
squeal_samples[27674]=52871;
squeal_samples[27675]=47324;
squeal_samples[27676]=41924;
squeal_samples[27677]=36879;
squeal_samples[27678]=32151;
squeal_samples[27679]=27726;
squeal_samples[27680]=23590;
squeal_samples[27681]=19715;
squeal_samples[27682]=16091;
squeal_samples[27683]=12695;
squeal_samples[27684]=9523;
squeal_samples[27685]=6556;
squeal_samples[27686]=4896;
squeal_samples[27687]=7509;
squeal_samples[27688]=10399;
squeal_samples[27689]=13170;
squeal_samples[27690]=15815;
squeal_samples[27691]=18353;
squeal_samples[27692]=20764;
squeal_samples[27693]=23084;
squeal_samples[27694]=25283;
squeal_samples[27695]=27410;
squeal_samples[27696]=29422;
squeal_samples[27697]=31352;
squeal_samples[27698]=33196;
squeal_samples[27699]=34953;
squeal_samples[27700]=36637;
squeal_samples[27701]=38241;
squeal_samples[27702]=39779;
squeal_samples[27703]=41241;
squeal_samples[27704]=42645;
squeal_samples[27705]=43976;
squeal_samples[27706]=45254;
squeal_samples[27707]=46474;
squeal_samples[27708]=47635;
squeal_samples[27709]=48750;
squeal_samples[27710]=49808;
squeal_samples[27711]=50823;
squeal_samples[27712]=51793;
squeal_samples[27713]=52720;
squeal_samples[27714]=53607;
squeal_samples[27715]=53972;
squeal_samples[27716]=49432;
squeal_samples[27717]=43897;
squeal_samples[27718]=38723;
squeal_samples[27719]=33879;
squeal_samples[27720]=29337;
squeal_samples[27721]=25098;
squeal_samples[27722]=21124;
squeal_samples[27723]=17406;
squeal_samples[27724]=13937;
squeal_samples[27725]=10676;
squeal_samples[27726]=7633;
squeal_samples[27727]=4967;
squeal_samples[27728]=6376;
squeal_samples[27729]=9318;
squeal_samples[27730]=12131;
squeal_samples[27731]=14827;
squeal_samples[27732]=17400;
squeal_samples[27733]=19866;
squeal_samples[27734]=22211;
squeal_samples[27735]=24462;
squeal_samples[27736]=26613;
squeal_samples[27737]=28664;
squeal_samples[27738]=30628;
squeal_samples[27739]=32502;
squeal_samples[27740]=34290;
squeal_samples[27741]=36001;
squeal_samples[27742]=37640;
squeal_samples[27743]=39195;
squeal_samples[27744]=40691;
squeal_samples[27745]=42108;
squeal_samples[27746]=43473;
squeal_samples[27747]=44770;
squeal_samples[27748]=46011;
squeal_samples[27749]=47198;
squeal_samples[27750]=48323;
squeal_samples[27751]=49406;
squeal_samples[27752]=50437;
squeal_samples[27753]=51429;
squeal_samples[27754]=52364;
squeal_samples[27755]=53271;
squeal_samples[27756]=54124;
squeal_samples[27757]=51593;
squeal_samples[27758]=45915;
squeal_samples[27759]=40616;
squeal_samples[27760]=35637;
squeal_samples[27761]=31000;
squeal_samples[27762]=26640;
squeal_samples[27763]=22576;
squeal_samples[27764]=18763;
squeal_samples[27765]=15199;
squeal_samples[27766]=11862;
squeal_samples[27767]=8742;
squeal_samples[27768]=5818;
squeal_samples[27769]=5279;
squeal_samples[27770]=8218;
squeal_samples[27771]=11082;
squeal_samples[27772]=13823;
squeal_samples[27773]=16437;
squeal_samples[27774]=18943;
squeal_samples[27775]=21331;
squeal_samples[27776]=23615;
squeal_samples[27777]=25804;
squeal_samples[27778]=27892;
squeal_samples[27779]=29891;
squeal_samples[27780]=31794;
squeal_samples[27781]=33619;
squeal_samples[27782]=35359;
squeal_samples[27783]=37020;
squeal_samples[27784]=38611;
squeal_samples[27785]=40123;
squeal_samples[27786]=41573;
squeal_samples[27787]=42957;
squeal_samples[27788]=44279;
squeal_samples[27789]=45541;
squeal_samples[27790]=46744;
squeal_samples[27791]=47895;
squeal_samples[27792]=48999;
squeal_samples[27793]=50044;
squeal_samples[27794]=51054;
squeal_samples[27795]=52006;
squeal_samples[27796]=52924;
squeal_samples[27797]=53799;
squeal_samples[27798]=53311;
squeal_samples[27799]=47990;
squeal_samples[27800]=42549;
squeal_samples[27801]=37457;
squeal_samples[27802]=32692;
squeal_samples[27803]=28231;
squeal_samples[27804]=24054;
squeal_samples[27805]=20154;
squeal_samples[27806]=16497;
squeal_samples[27807]=13072;
squeal_samples[27808]=9877;
squeal_samples[27809]=6878;
squeal_samples[27810]=4799;
squeal_samples[27811]=7102;
squeal_samples[27812]=10014;
squeal_samples[27813]=12793;
squeal_samples[27814]=15455;
squeal_samples[27815]=18003;
squeal_samples[27816]=20438;
squeal_samples[27817]=22760;
squeal_samples[27818]=24981;
squeal_samples[27819]=27112;
squeal_samples[27820]=29140;
squeal_samples[27821]=31083;
squeal_samples[27822]=32934;
squeal_samples[27823]=34704;
squeal_samples[27824]=36393;
squeal_samples[27825]=38015;
squeal_samples[27826]=39551;
squeal_samples[27827]=41031;
squeal_samples[27828]=42435;
squeal_samples[27829]=43780;
squeal_samples[27830]=45062;
squeal_samples[27831]=46287;
squeal_samples[27832]=47462;
squeal_samples[27833]=48576;
squeal_samples[27834]=49647;
squeal_samples[27835]=50661;
squeal_samples[27836]=51646;
squeal_samples[27837]=52571;
squeal_samples[27838]=53462;
squeal_samples[27839]=54264;
squeal_samples[27840]=50935;
squeal_samples[27841]=45302;
squeal_samples[27842]=40038;
squeal_samples[27843]=35100;
squeal_samples[27844]=30491;
squeal_samples[27845]=26164;
squeal_samples[27846]=22126;
squeal_samples[27847]=18347;
squeal_samples[27848]=14804;
squeal_samples[27849]=11495;
squeal_samples[27850]=8388;
squeal_samples[27851]=5496;
squeal_samples[27852]=5631;
squeal_samples[27853]=8606;
squeal_samples[27854]=11446;
squeal_samples[27855]=14166;
squeal_samples[27856]=16771;
squeal_samples[27857]=19259;
squeal_samples[27858]=21633;
squeal_samples[27859]=23910;
squeal_samples[27860]=26076;
squeal_samples[27861]=28162;
squeal_samples[27862]=30133;
squeal_samples[27863]=32037;
squeal_samples[27864]=33841;
squeal_samples[27865]=35579;
squeal_samples[27866]=37222;
squeal_samples[27867]=38806;
squeal_samples[27868]=40306;
squeal_samples[27869]=41752;
squeal_samples[27870]=43122;
squeal_samples[27871]=44437;
squeal_samples[27872]=45690;
squeal_samples[27873]=46884;
squeal_samples[27874]=48032;
squeal_samples[27875]=49119;
squeal_samples[27876]=50165;
squeal_samples[27877]=51164;
squeal_samples[27878]=52116;
squeal_samples[27879]=53023;
squeal_samples[27880]=53899;
squeal_samples[27881]=53399;
squeal_samples[27882]=48071;
squeal_samples[27883]=42625;
squeal_samples[27884]=37524;
squeal_samples[27885]=32758;
squeal_samples[27886]=28288;
squeal_samples[27887]=24107;
squeal_samples[27888]=20203;
squeal_samples[27889]=16537;
squeal_samples[27890]=13116;
squeal_samples[27891]=9913;
squeal_samples[27892]=6909;
squeal_samples[27893]=4831;
squeal_samples[27894]=7128;
squeal_samples[27895]=10040;
squeal_samples[27896]=12818;
squeal_samples[27897]=15477;
squeal_samples[27898]=18021;
squeal_samples[27899]=20457;
squeal_samples[27900]=22771;
squeal_samples[27901]=24999;
squeal_samples[27902]=27121;
squeal_samples[27903]=29149;
squeal_samples[27904]=31089;
squeal_samples[27905]=32942;
squeal_samples[27906]=34713;
squeal_samples[27907]=36400;
squeal_samples[27908]=38016;
squeal_samples[27909]=39559;
squeal_samples[27910]=41027;
squeal_samples[27911]=42434;
squeal_samples[27912]=43780;
squeal_samples[27913]=45059;
squeal_samples[27914]=46288;
squeal_samples[27915]=47452;
squeal_samples[27916]=48575;
squeal_samples[27917]=49639;
squeal_samples[27918]=50661;
squeal_samples[27919]=51628;
squeal_samples[27920]=52569;
squeal_samples[27921]=53454;
squeal_samples[27922]=54251;
squeal_samples[27923]=50925;
squeal_samples[27924]=45288;
squeal_samples[27925]=40028;
squeal_samples[27926]=35088;
squeal_samples[27927]=30478;
squeal_samples[27928]=26152;
squeal_samples[27929]=22110;
squeal_samples[27930]=18327;
squeal_samples[27931]=14791;
squeal_samples[27932]=11472;
squeal_samples[27933]=8377;
squeal_samples[27934]=5471;
squeal_samples[27935]=5621;
squeal_samples[27936]=8584;
squeal_samples[27937]=11430;
squeal_samples[27938]=14150;
squeal_samples[27939]=16751;
squeal_samples[27940]=19243;
squeal_samples[27941]=21618;
squeal_samples[27942]=23883;
squeal_samples[27943]=26064;
squeal_samples[27944]=28133;
squeal_samples[27945]=30122;
squeal_samples[27946]=32015;
squeal_samples[27947]=33826;
squeal_samples[27948]=35555;
squeal_samples[27949]=37206;
squeal_samples[27950]=38783;
squeal_samples[27951]=40289;
squeal_samples[27952]=41728;
squeal_samples[27953]=43100;
squeal_samples[27954]=44414;
squeal_samples[27955]=45669;
squeal_samples[27956]=46865;
squeal_samples[27957]=48009;
squeal_samples[27958]=49102;
squeal_samples[27959]=50148;
squeal_samples[27960]=51141;
squeal_samples[27961]=52093;
squeal_samples[27962]=53001;
squeal_samples[27963]=53874;
squeal_samples[27964]=53385;
squeal_samples[27965]=48050;
squeal_samples[27966]=42605;
squeal_samples[27967]=37505;
squeal_samples[27968]=32737;
squeal_samples[27969]=28264;
squeal_samples[27970]=24085;
squeal_samples[27971]=20180;
squeal_samples[27972]=16520;
squeal_samples[27973]=13093;
squeal_samples[27974]=9889;
squeal_samples[27975]=6890;
squeal_samples[27976]=4804;
squeal_samples[27977]=7110;
squeal_samples[27978]=10012;
squeal_samples[27979]=12800;
squeal_samples[27980]=15450;
squeal_samples[27981]=18004;
squeal_samples[27982]=20427;
squeal_samples[27983]=22755;
squeal_samples[27984]=24972;
squeal_samples[27985]=27101;
squeal_samples[27986]=29124;
squeal_samples[27987]=31067;
squeal_samples[27988]=32919;
squeal_samples[27989]=34691;
squeal_samples[27990]=36377;
squeal_samples[27991]=37994;
squeal_samples[27992]=39534;
squeal_samples[27993]=41007;
squeal_samples[27994]=42410;
squeal_samples[27995]=43756;
squeal_samples[27996]=45040;
squeal_samples[27997]=46262;
squeal_samples[27998]=47431;
squeal_samples[27999]=48552;
squeal_samples[28000]=49616;
squeal_samples[28001]=50639;
squeal_samples[28002]=51610;
squeal_samples[28003]=52547;
squeal_samples[28004]=53429;
squeal_samples[28005]=54233;
squeal_samples[28006]=50896;
squeal_samples[28007]=45271;
squeal_samples[28008]=40000;
squeal_samples[28009]=35070;
squeal_samples[28010]=30453;
squeal_samples[28011]=26130;
squeal_samples[28012]=22087;
squeal_samples[28013]=18303;
squeal_samples[28014]=14771;
squeal_samples[28015]=11448;
squeal_samples[28016]=8354;
squeal_samples[28017]=5451;
squeal_samples[28018]=5594;
squeal_samples[28019]=8565;
squeal_samples[28020]=11405;
squeal_samples[28021]=14128;
squeal_samples[28022]=16729;
squeal_samples[28023]=19220;
squeal_samples[28024]=21595;
squeal_samples[28025]=23861;
squeal_samples[28026]=26039;
squeal_samples[28027]=28114;
squeal_samples[28028]=30095;
squeal_samples[28029]=31996;
squeal_samples[28030]=33802;
squeal_samples[28031]=35531;
squeal_samples[28032]=37186;
squeal_samples[28033]=38758;
squeal_samples[28034]=40266;
squeal_samples[28035]=41708;
squeal_samples[28036]=43075;
squeal_samples[28037]=44393;
squeal_samples[28038]=45643;
squeal_samples[28039]=46846;
squeal_samples[28040]=47984;
squeal_samples[28041]=49082;
squeal_samples[28042]=50123;
squeal_samples[28043]=51119;
squeal_samples[28044]=52070;
squeal_samples[28045]=52980;
squeal_samples[28046]=53851;
squeal_samples[28047]=53361;
squeal_samples[28048]=48030;
squeal_samples[28049]=42578;
squeal_samples[28050]=37489;
squeal_samples[28051]=32708;
squeal_samples[28052]=28246;
squeal_samples[28053]=24059;
squeal_samples[28054]=20158;
squeal_samples[28055]=16499;
squeal_samples[28056]=13069;
squeal_samples[28057]=9867;
squeal_samples[28058]=6867;
squeal_samples[28059]=4781;
squeal_samples[28060]=7087;
squeal_samples[28061]=9990;
squeal_samples[28062]=12777;
squeal_samples[28063]=15429;
squeal_samples[28064]=17978;
squeal_samples[28065]=20409;
squeal_samples[28066]=22728;
squeal_samples[28067]=24952;
squeal_samples[28068]=27076;
squeal_samples[28069]=29104;
squeal_samples[28070]=31043;
squeal_samples[28071]=32899;
squeal_samples[28072]=34665;
squeal_samples[28073]=36356;
squeal_samples[28074]=37971;
squeal_samples[28075]=39511;
squeal_samples[28076]=40986;
squeal_samples[28077]=42385;
squeal_samples[28078]=43738;
squeal_samples[28079]=45010;
squeal_samples[28080]=46246;
squeal_samples[28081]=47405;
squeal_samples[28082]=48529;
squeal_samples[28083]=49596;
squeal_samples[28084]=50613;
squeal_samples[28085]=51590;
squeal_samples[28086]=52523;
squeal_samples[28087]=53407;
squeal_samples[28088]=54209;
squeal_samples[28089]=50875;
squeal_samples[28090]=45249;
squeal_samples[28091]=39975;
squeal_samples[28092]=35050;
squeal_samples[28093]=30426;
squeal_samples[28094]=26113;
squeal_samples[28095]=22059;
squeal_samples[28096]=18286;
squeal_samples[28097]=14744;
squeal_samples[28098]=11426;
squeal_samples[28099]=8332;
squeal_samples[28100]=5427;
squeal_samples[28101]=5573;
squeal_samples[28102]=8542;
squeal_samples[28103]=11382;
squeal_samples[28104]=14105;
squeal_samples[28105]=16706;
squeal_samples[28106]=19199;
squeal_samples[28107]=21570;
squeal_samples[28108]=23841;
squeal_samples[28109]=26015;
squeal_samples[28110]=28090;
squeal_samples[28111]=30076;
squeal_samples[28112]=31969;
squeal_samples[28113]=33783;
squeal_samples[28114]=35507;
squeal_samples[28115]=37163;
squeal_samples[28116]=38735;
squeal_samples[28117]=40246;
squeal_samples[28118]=41680;
squeal_samples[28119]=43058;
squeal_samples[28120]=44366;
squeal_samples[28121]=45624;
squeal_samples[28122]=46821;
squeal_samples[28123]=47962;
squeal_samples[28124]=49059;
squeal_samples[28125]=50100;
squeal_samples[28126]=51098;
squeal_samples[28127]=52046;
squeal_samples[28128]=52957;
squeal_samples[28129]=53829;
squeal_samples[28130]=53338;
squeal_samples[28131]=48008;
squeal_samples[28132]=42555;
squeal_samples[28133]=37464;
squeal_samples[28134]=32689;
squeal_samples[28135]=28220;
squeal_samples[28136]=24040;
squeal_samples[28137]=20133;
squeal_samples[28138]=16475;
squeal_samples[28139]=13050;
squeal_samples[28140]=9841;
squeal_samples[28141]=6846;
squeal_samples[28142]=4758;
squeal_samples[28143]=7064;
squeal_samples[28144]=9968;
squeal_samples[28145]=12754;
squeal_samples[28146]=15405;
squeal_samples[28147]=17957;
squeal_samples[28148]=20386;
squeal_samples[28149]=22704;
squeal_samples[28150]=24932;
squeal_samples[28151]=27049;
squeal_samples[28152]=29086;
squeal_samples[28153]=31017;
squeal_samples[28154]=32877;
squeal_samples[28155]=34642;
squeal_samples[28156]=36334;
squeal_samples[28157]=37946;
squeal_samples[28158]=39493;
squeal_samples[28159]=40957;
squeal_samples[28160]=42367;
squeal_samples[28161]=43712;
squeal_samples[28162]=44990;
squeal_samples[28163]=46221;
squeal_samples[28164]=47383;
squeal_samples[28165]=48506;
squeal_samples[28166]=49573;
squeal_samples[28167]=50590;
squeal_samples[28168]=51568;
squeal_samples[28169]=52498;
squeal_samples[28170]=53386;
squeal_samples[28171]=54238;
squeal_samples[28172]=51684;
squeal_samples[28173]=46003;
squeal_samples[28174]=40681;
squeal_samples[28175]=35703;
squeal_samples[28176]=31044;
squeal_samples[28177]=26681;
squeal_samples[28178]=22601;
squeal_samples[28179]=18781;
squeal_samples[28180]=15209;
squeal_samples[28181]=11864;
squeal_samples[28182]=8735;
squeal_samples[28183]=5802;
squeal_samples[28184]=5264;
squeal_samples[28185]=8193;
squeal_samples[28186]=11061;
squeal_samples[28187]=13785;
squeal_samples[28188]=16409;
squeal_samples[28189]=18902;
squeal_samples[28190]=21289;
squeal_samples[28191]=23571;
squeal_samples[28192]=25757;
squeal_samples[28193]=27842;
squeal_samples[28194]=29837;
squeal_samples[28195]=31741;
squeal_samples[28196]=33556;
squeal_samples[28197]=35304;
squeal_samples[28198]=36958;
squeal_samples[28199]=38546;
squeal_samples[28200]=40059;
squeal_samples[28201]=41501;
squeal_samples[28202]=42887;
squeal_samples[28203]=44205;
squeal_samples[28204]=45463;
squeal_samples[28205]=46668;
squeal_samples[28206]=47822;
squeal_samples[28207]=48912;
squeal_samples[28208]=49968;
squeal_samples[28209]=50963;
squeal_samples[28210]=51919;
squeal_samples[28211]=52840;
squeal_samples[28212]=53706;
squeal_samples[28213]=54076;
squeal_samples[28214]=49502;
squeal_samples[28215]=43964;
squeal_samples[28216]=38776;
squeal_samples[28217]=33914;
squeal_samples[28218]=29372;
squeal_samples[28219]=25111;
squeal_samples[28220]=21135;
squeal_samples[28221]=17405;
squeal_samples[28222]=13923;
squeal_samples[28223]=10662;
squeal_samples[28224]=7609;
squeal_samples[28225]=4934;
squeal_samples[28226]=6342;
squeal_samples[28227]=9279;
squeal_samples[28228]=12087;
squeal_samples[28229]=14778;
squeal_samples[28230]=17345;
squeal_samples[28231]=19804;
squeal_samples[28232]=22151;
squeal_samples[28233]=24396;
squeal_samples[28234]=26542;
squeal_samples[28235]=28593;
squeal_samples[28236]=30551;
squeal_samples[28237]=32424;
squeal_samples[28238]=34215;
squeal_samples[28239]=35923;
squeal_samples[28240]=37553;
squeal_samples[28241]=39112;
squeal_samples[28242]=40604;
squeal_samples[28243]=42019;
squeal_samples[28244]=43383;
squeal_samples[28245]=44674;
squeal_samples[28246]=45914;
squeal_samples[28247]=47098;
squeal_samples[28248]=48224;
squeal_samples[28249]=49309;
squeal_samples[28250]=50331;
squeal_samples[28251]=51320;
squeal_samples[28252]=52255;
squeal_samples[28253]=53158;
squeal_samples[28254]=54017;
squeal_samples[28255]=52934;
squeal_samples[28256]=47377;
squeal_samples[28257]=41967;
squeal_samples[28258]=36908;
squeal_samples[28259]=32166;
squeal_samples[28260]=27729;
squeal_samples[28261]=23583;
squeal_samples[28262]=19697;
squeal_samples[28263]=16067;
squeal_samples[28264]=12661;
squeal_samples[28265]=9483;
squeal_samples[28266]=6504;
squeal_samples[28267]=4842;
squeal_samples[28268]=7444;
squeal_samples[28269]=10341;
squeal_samples[28270]=13096;
squeal_samples[28271]=15743;
squeal_samples[28272]=18274;
squeal_samples[28273]=20688;
squeal_samples[28274]=22997;
squeal_samples[28275]=25201;
squeal_samples[28276]=27309;
squeal_samples[28277]=29334;
squeal_samples[28278]=31253;
squeal_samples[28279]=33099;
squeal_samples[28280]=34853;
squeal_samples[28281]=36531;
squeal_samples[28282]=38138;
squeal_samples[28283]=39666;
squeal_samples[28284]=41134;
squeal_samples[28285]=42525;
squeal_samples[28286]=43863;
squeal_samples[28287]=45137;
squeal_samples[28288]=46352;
squeal_samples[28289]=47516;
squeal_samples[28290]=48625;
squeal_samples[28291]=49689;
squeal_samples[28292]=50695;
squeal_samples[28293]=51667;
squeal_samples[28294]=52586;
squeal_samples[28295]=53476;
squeal_samples[28296]=54264;
squeal_samples[28297]=50934;
squeal_samples[28298]=45289;
squeal_samples[28299]=40021;
squeal_samples[28300]=35082;
squeal_samples[28301]=30453;
squeal_samples[28302]=26135;
squeal_samples[28303]=22082;
squeal_samples[28304]=18296;
squeal_samples[28305]=14754;
squeal_samples[28306]=11429;
squeal_samples[28307]=8335;
squeal_samples[28308]=5424;
squeal_samples[28309]=5567;
squeal_samples[28310]=8531;
squeal_samples[28311]=11377;
squeal_samples[28312]=14090;
squeal_samples[28313]=16694;
squeal_samples[28314]=19178;
squeal_samples[28315]=21554;
squeal_samples[28316]=23819;
squeal_samples[28317]=25994;
squeal_samples[28318]=28064;
squeal_samples[28319]=30052;
squeal_samples[28320]=31946;
squeal_samples[28321]=33751;
squeal_samples[28322]=35480;
squeal_samples[28323]=37125;
squeal_samples[28324]=38709;
squeal_samples[28325]=40207;
squeal_samples[28326]=41650;
squeal_samples[28327]=43023;
squeal_samples[28328]=44336;
squeal_samples[28329]=45585;
squeal_samples[28330]=46782;
squeal_samples[28331]=47927;
squeal_samples[28332]=49018;
squeal_samples[28333]=50061;
squeal_samples[28334]=51056;
squeal_samples[28335]=52005;
squeal_samples[28336]=52917;
squeal_samples[28337]=53781;
squeal_samples[28338]=53767;
squeal_samples[28339]=48758;
squeal_samples[28340]=43263;
squeal_samples[28341]=38115;
squeal_samples[28342]=33302;
squeal_samples[28343]=28786;
squeal_samples[28344]=24570;
squeal_samples[28345]=20626;
squeal_samples[28346]=16929;
squeal_samples[28347]=13469;
squeal_samples[28348]=10232;
squeal_samples[28349]=7206;
squeal_samples[28350]=4779;
squeal_samples[28351]=6685;
squeal_samples[28352]=9602;
squeal_samples[28353]=12398;
squeal_samples[28354]=15068;
squeal_samples[28355]=17626;
squeal_samples[28356]=20076;
squeal_samples[28357]=22402;
squeal_samples[28358]=24636;
squeal_samples[28359]=26773;
squeal_samples[28360]=28808;
squeal_samples[28361]=30757;
squeal_samples[28362]=32618;
squeal_samples[28363]=34397;
squeal_samples[28364]=36096;
squeal_samples[28365]=37720;
squeal_samples[28366]=39269;
squeal_samples[28367]=40747;
squeal_samples[28368]=42162;
squeal_samples[28369]=43507;
squeal_samples[28370]=44802;
squeal_samples[28371]=46030;
squeal_samples[28372]=47206;
squeal_samples[28373]=48326;
squeal_samples[28374]=49404;
squeal_samples[28375]=50424;
squeal_samples[28376]=51404;
squeal_samples[28377]=52337;
squeal_samples[28378]=53237;
squeal_samples[28379]=54088;
squeal_samples[28380]=52324;
squeal_samples[28381]=46647;
squeal_samples[28382]=41281;
squeal_samples[28383]=36263;
squeal_samples[28384]=31558;
squeal_samples[28385]=27168;
squeal_samples[28386]=23043;
squeal_samples[28387]=19203;
squeal_samples[28388]=15589;
squeal_samples[28389]=12222;
squeal_samples[28390]=9061;
squeal_samples[28391]=6115;
squeal_samples[28392]=4961;
squeal_samples[28393]=7787;
squeal_samples[28394]=10647;
squeal_samples[28395]=13405;
squeal_samples[28396]=16027;
squeal_samples[28397]=18543;
squeal_samples[28398]=20945;
squeal_samples[28399]=23238;
squeal_samples[28400]=25438;
squeal_samples[28401]=27539;
squeal_samples[28402]=29538;
squeal_samples[28403]=31459;
squeal_samples[28404]=33284;
squeal_samples[28405]=35031;
squeal_samples[28406]=36706;
squeal_samples[28407]=38295;
squeal_samples[28408]=39822;
squeal_samples[28409]=41269;
squeal_samples[28410]=42664;
squeal_samples[28411]=43988;
squeal_samples[28412]=45258;
squeal_samples[28413]=46462;
squeal_samples[28414]=47625;
squeal_samples[28415]=48723;
squeal_samples[28416]=49783;
squeal_samples[28417]=50788;
squeal_samples[28418]=51750;
squeal_samples[28419]=52670;
squeal_samples[28420]=53547;
squeal_samples[28421]=54176;
squeal_samples[28422]=50172;
squeal_samples[28423]=44581;
squeal_samples[28424]=39348;
squeal_samples[28425]=34453;
squeal_samples[28426]=29864;
squeal_samples[28427]=25581;
squeal_samples[28428]=21558;
squeal_samples[28429]=17807;
squeal_samples[28430]=14291;
squeal_samples[28431]=10999;
squeal_samples[28432]=7926;
squeal_samples[28433]=5086;
squeal_samples[28434]=5912;
squeal_samples[28435]=8863;
squeal_samples[28436]=11691;
squeal_samples[28437]=14386;
squeal_samples[28438]=16983;
squeal_samples[28439]=19446;
squeal_samples[28440]=21808;
squeal_samples[28441]=24064;
squeal_samples[28442]=26224;
squeal_samples[28443]=28286;
squeal_samples[28444]=30257;
squeal_samples[28445]=32140;
squeal_samples[28446]=33940;
squeal_samples[28447]=35657;
squeal_samples[28448]=37299;
squeal_samples[28449]=38862;
squeal_samples[28450]=40362;
squeal_samples[28451]=41791;
squeal_samples[28452]=43155;
squeal_samples[28453]=44463;
squeal_samples[28454]=45703;
squeal_samples[28455]=46898;
squeal_samples[28456]=48024;
squeal_samples[28457]=49118;
squeal_samples[28458]=50150;
squeal_samples[28459]=51142;
squeal_samples[28460]=52086;
squeal_samples[28461]=52992;
squeal_samples[28462]=53856;
squeal_samples[28463]=53359;
squeal_samples[28464]=48016;
squeal_samples[28465]=42572;
squeal_samples[28466]=37462;
squeal_samples[28467]=32688;
squeal_samples[28468]=28209;
squeal_samples[28469]=24026;
squeal_samples[28470]=20113;
squeal_samples[28471]=16450;
squeal_samples[28472]=13017;
squeal_samples[28473]=9813;
squeal_samples[28474]=6807;
squeal_samples[28475]=4719;
squeal_samples[28476]=7021;
squeal_samples[28477]=9921;
squeal_samples[28478]=12706;
squeal_samples[28479]=15360;
squeal_samples[28480]=17908;
squeal_samples[28481]=20334;
squeal_samples[28482]=22652;
squeal_samples[28483]=24877;
squeal_samples[28484]=27002;
squeal_samples[28485]=29022;
squeal_samples[28486]=30963;
squeal_samples[28487]=32811;
squeal_samples[28488]=34581;
squeal_samples[28489]=36269;
squeal_samples[28490]=37880;
squeal_samples[28491]=39420;
squeal_samples[28492]=40892;
squeal_samples[28493]=42296;
squeal_samples[28494]=43643;
squeal_samples[28495]=44922;
squeal_samples[28496]=46147;
squeal_samples[28497]=47313;
squeal_samples[28498]=48433;
squeal_samples[28499]=49497;
squeal_samples[28500]=50516;
squeal_samples[28501]=51489;
squeal_samples[28502]=52417;
squeal_samples[28503]=53312;
squeal_samples[28504]=54156;
squeal_samples[28505]=52389;
squeal_samples[28506]=46704;
squeal_samples[28507]=41336;
squeal_samples[28508]=36306;
squeal_samples[28509]=31605;
squeal_samples[28510]=27199;
squeal_samples[28511]=23081;
squeal_samples[28512]=19222;
squeal_samples[28513]=15619;
squeal_samples[28514]=12240;
squeal_samples[28515]=9077;
squeal_samples[28516]=6129;
squeal_samples[28517]=4972;
squeal_samples[28518]=7794;
squeal_samples[28519]=10659;
squeal_samples[28520]=13413;
squeal_samples[28521]=16030;
squeal_samples[28522]=18551;
squeal_samples[28523]=20939;
squeal_samples[28524]=23239;
squeal_samples[28525]=25437;
squeal_samples[28526]=27530;
squeal_samples[28527]=29534;
squeal_samples[28528]=31451;
squeal_samples[28529]=33275;
squeal_samples[28530]=35028;
squeal_samples[28531]=36689;
squeal_samples[28532]=38288;
squeal_samples[28533]=39805;
squeal_samples[28534]=41260;
squeal_samples[28535]=42648;
squeal_samples[28536]=43973;
squeal_samples[28537]=45245;
squeal_samples[28538]=46444;
squeal_samples[28539]=47608;
squeal_samples[28540]=48703;
squeal_samples[28541]=49762;
squeal_samples[28542]=50768;
squeal_samples[28543]=51729;
squeal_samples[28544]=52644;
squeal_samples[28545]=53531;
squeal_samples[28546]=54314;
squeal_samples[28547]=50970;
squeal_samples[28548]=45328;
squeal_samples[28549]=40044;
squeal_samples[28550]=35099;
squeal_samples[28551]=30476;
squeal_samples[28552]=26139;
squeal_samples[28553]=22088;
squeal_samples[28554]=18291;
squeal_samples[28555]=14752;
squeal_samples[28556]=11422;
squeal_samples[28557]=8319;
squeal_samples[28558]=5408;
squeal_samples[28559]=5545;
squeal_samples[28560]=8515;
squeal_samples[28561]=11350;
squeal_samples[28562]=14067;
squeal_samples[28563]=16669;
squeal_samples[28564]=19149;
squeal_samples[28565]=21523;
squeal_samples[28566]=23791;
squeal_samples[28567]=25961;
squeal_samples[28568]=28037;
squeal_samples[28569]=30010;
squeal_samples[28570]=31905;
squeal_samples[28571]=33712;
squeal_samples[28572]=35437;
squeal_samples[28573]=37086;
squeal_samples[28574]=38667;
squeal_samples[28575]=40167;
squeal_samples[28576]=41609;
squeal_samples[28577]=42977;
squeal_samples[28578]=44289;
squeal_samples[28579]=45540;
squeal_samples[28580]=46735;
squeal_samples[28581]=47876;
squeal_samples[28582]=48965;
squeal_samples[28583]=50010;
squeal_samples[28584]=51003;
squeal_samples[28585]=51954;
squeal_samples[28586]=52866;
squeal_samples[28587]=53728;
squeal_samples[28588]=54084;
squeal_samples[28589]=49511;
squeal_samples[28590]=43964;
squeal_samples[28591]=38767;
squeal_samples[28592]=33907;
squeal_samples[28593]=29347;
squeal_samples[28594]=25095;
squeal_samples[28595]=21100;
squeal_samples[28596]=17377;
squeal_samples[28597]=13886;
squeal_samples[28598]=10619;
squeal_samples[28599]=7561;
squeal_samples[28600]=4882;
squeal_samples[28601]=6288;
squeal_samples[28602]=9229;
squeal_samples[28603]=12026;
squeal_samples[28604]=14722;
squeal_samples[28605]=17283;
squeal_samples[28606]=19750;
squeal_samples[28607]=22085;
squeal_samples[28608]=24333;
squeal_samples[28609]=26478;
squeal_samples[28610]=28524;
squeal_samples[28611]=30481;
squeal_samples[28612]=32357;
squeal_samples[28613]=34138;
squeal_samples[28614]=35850;
squeal_samples[28615]=37476;
squeal_samples[28616]=39036;
squeal_samples[28617]=40519;
squeal_samples[28618]=41945;
squeal_samples[28619]=43297;
squeal_samples[28620]=44598;
squeal_samples[28621]=45832;
squeal_samples[28622]=47012;
squeal_samples[28623]=48142;
squeal_samples[28624]=49219;
squeal_samples[28625]=50250;
squeal_samples[28626]=51230;
squeal_samples[28627]=52172;
squeal_samples[28628]=53071;
squeal_samples[28629]=53932;
squeal_samples[28630]=53424;
squeal_samples[28631]=48083;
squeal_samples[28632]=42622;
squeal_samples[28633]=37512;
squeal_samples[28634]=32726;
squeal_samples[28635]=28248;
squeal_samples[28636]=24054;
squeal_samples[28637]=20141;
squeal_samples[28638]=16469;
squeal_samples[28639]=13037;
squeal_samples[28640]=9822;
squeal_samples[28641]=6816;
squeal_samples[28642]=4727;
squeal_samples[28643]=7026;
squeal_samples[28644]=9924;
squeal_samples[28645]=12705;
squeal_samples[28646]=15358;
squeal_samples[28647]=17899;
squeal_samples[28648]=20334;
squeal_samples[28649]=22645;
squeal_samples[28650]=24864;
squeal_samples[28651]=26989;
squeal_samples[28652]=29010;
squeal_samples[28653]=30948;
squeal_samples[28654]=32803;
squeal_samples[28655]=34559;
squeal_samples[28656]=36253;
squeal_samples[28657]=37860;
squeal_samples[28658]=39403;
squeal_samples[28659]=40874;
squeal_samples[28660]=42278;
squeal_samples[28661]=43620;
squeal_samples[28662]=44897;
squeal_samples[28663]=46125;
squeal_samples[28664]=47284;
squeal_samples[28665]=48409;
squeal_samples[28666]=49469;
squeal_samples[28667]=50487;
squeal_samples[28668]=51460;
squeal_samples[28669]=52388;
squeal_samples[28670]=53279;
squeal_samples[28671]=54126;
squeal_samples[28672]=52356;
squeal_samples[28673]=46667;
squeal_samples[28674]=41305;
squeal_samples[28675]=36269;
squeal_samples[28676]=31574;
squeal_samples[28677]=27162;
squeal_samples[28678]=23042;
squeal_samples[28679]=19188;
squeal_samples[28680]=15580;
squeal_samples[28681]=12198;
squeal_samples[28682]=9046;
squeal_samples[28683]=6086;
squeal_samples[28684]=4936;
squeal_samples[28685]=7751;
squeal_samples[28686]=10622;
squeal_samples[28687]=13365;
squeal_samples[28688]=15994;
squeal_samples[28689]=18508;
squeal_samples[28690]=20902;
squeal_samples[28691]=23198;
squeal_samples[28692]=25392;
squeal_samples[28693]=27491;
squeal_samples[28694]=29494;
squeal_samples[28695]=31411;
squeal_samples[28696]=33231;
squeal_samples[28697]=34982;
squeal_samples[28698]=36651;
squeal_samples[28699]=38241;
squeal_samples[28700]=39766;
squeal_samples[28701]=41221;
squeal_samples[28702]=42602;
squeal_samples[28703]=43936;
squeal_samples[28704]=45196;
squeal_samples[28705]=46408;
squeal_samples[28706]=47566;
squeal_samples[28707]=48664;
squeal_samples[28708]=49722;
squeal_samples[28709]=50725;
squeal_samples[28710]=51686;
squeal_samples[28711]=52608;
squeal_samples[28712]=53483;
squeal_samples[28713]=54270;
squeal_samples[28714]=50931;
squeal_samples[28715]=45282;
squeal_samples[28716]=40004;
squeal_samples[28717]=35056;
squeal_samples[28718]=30429;
squeal_samples[28719]=26095;
squeal_samples[28720]=22042;
squeal_samples[28721]=18252;
squeal_samples[28722]=14707;
squeal_samples[28723]=11377;
squeal_samples[28724]=8274;
squeal_samples[28725]=5363;
squeal_samples[28726]=5500;
squeal_samples[28727]=8469;
squeal_samples[28728]=11307;
squeal_samples[28729]=14021;
squeal_samples[28730]=16623;
squeal_samples[28731]=19106;
squeal_samples[28732]=21476;
squeal_samples[28733]=23748;
squeal_samples[28734]=25915;
squeal_samples[28735]=27992;
squeal_samples[28736]=29970;
squeal_samples[28737]=31862;
squeal_samples[28738]=33664;
squeal_samples[28739]=35395;
squeal_samples[28740]=37039;
squeal_samples[28741]=38623;
squeal_samples[28742]=40122;
squeal_samples[28743]=41563;
squeal_samples[28744]=42933;
squeal_samples[28745]=44244;
squeal_samples[28746]=45494;
squeal_samples[28747]=46692;
squeal_samples[28748]=47827;
squeal_samples[28749]=48925;
squeal_samples[28750]=49961;
squeal_samples[28751]=50961;
squeal_samples[28752]=51908;
squeal_samples[28753]=52820;
squeal_samples[28754]=53684;
squeal_samples[28755]=54040;
squeal_samples[28756]=49463;
squeal_samples[28757]=43925;
squeal_samples[28758]=38716;
squeal_samples[28759]=33865;
squeal_samples[28760]=29302;
squeal_samples[28761]=25049;
squeal_samples[28762]=21057;
squeal_samples[28763]=17331;
squeal_samples[28764]=13840;
squeal_samples[28765]=10575;
squeal_samples[28766]=7517;
squeal_samples[28767]=4835;
squeal_samples[28768]=6246;
squeal_samples[28769]=9179;
squeal_samples[28770]=11988;
squeal_samples[28771]=14669;
squeal_samples[28772]=17246;
squeal_samples[28773]=19698;
squeal_samples[28774]=22044;
squeal_samples[28775]=24287;
squeal_samples[28776]=26433;
squeal_samples[28777]=28479;
squeal_samples[28778]=30436;
squeal_samples[28779]=32313;
squeal_samples[28780]=34091;
squeal_samples[28781]=35808;
squeal_samples[28782]=37428;
squeal_samples[28783]=38993;
squeal_samples[28784]=40473;
squeal_samples[28785]=41901;
squeal_samples[28786]=43252;
squeal_samples[28787]=44552;
squeal_samples[28788]=45788;
squeal_samples[28789]=46966;
squeal_samples[28790]=48097;
squeal_samples[28791]=49176;
squeal_samples[28792]=50203;
squeal_samples[28793]=51186;
squeal_samples[28794]=52127;
squeal_samples[28795]=53025;
squeal_samples[28796]=53888;
squeal_samples[28797]=53378;
squeal_samples[28798]=48041;
squeal_samples[28799]=42573;
squeal_samples[28800]=37470;
squeal_samples[28801]=32679;
squeal_samples[28802]=28204;
squeal_samples[28803]=24010;
squeal_samples[28804]=20094;
squeal_samples[28805]=16425;
squeal_samples[28806]=12993;
squeal_samples[28807]=9774;
squeal_samples[28808]=6776;
squeal_samples[28809]=4676;
squeal_samples[28810]=6987;
squeal_samples[28811]=9874;
squeal_samples[28812]=12664;
squeal_samples[28813]=15309;
squeal_samples[28814]=17858;
squeal_samples[28815]=20286;
squeal_samples[28816]=22601;
squeal_samples[28817]=24820;
squeal_samples[28818]=26942;
squeal_samples[28819]=28966;
squeal_samples[28820]=30905;
squeal_samples[28821]=32753;
squeal_samples[28822]=34519;
squeal_samples[28823]=36204;
squeal_samples[28824]=37818;
squeal_samples[28825]=39357;
squeal_samples[28826]=40828;
squeal_samples[28827]=42234;
squeal_samples[28828]=43573;
squeal_samples[28829]=44856;
squeal_samples[28830]=46074;
squeal_samples[28831]=47244;
squeal_samples[28832]=48361;
squeal_samples[28833]=49424;
squeal_samples[28834]=50443;
squeal_samples[28835]=51413;
squeal_samples[28836]=52344;
squeal_samples[28837]=53232;
squeal_samples[28838]=54082;
squeal_samples[28839]=52987;
squeal_samples[28840]=47415;
squeal_samples[28841]=41992;
squeal_samples[28842]=36921;
squeal_samples[28843]=32166;
squeal_samples[28844]=27729;
squeal_samples[28845]=23559;
squeal_samples[28846]=19681;
squeal_samples[28847]=16030;
squeal_samples[28848]=12623;
squeal_samples[28849]=9434;
squeal_samples[28850]=6444;
squeal_samples[28851]=4780;
squeal_samples[28852]=7382;
squeal_samples[28853]=10265;
squeal_samples[28854]=13028;
squeal_samples[28855]=15666;
squeal_samples[28856]=18191;
squeal_samples[28857]=20602;
squeal_samples[28858]=22904;
squeal_samples[28859]=25111;
squeal_samples[28860]=27221;
squeal_samples[28861]=29230;
squeal_samples[28862]=31154;
squeal_samples[28863]=32993;
squeal_samples[28864]=34743;
squeal_samples[28865]=36424;
squeal_samples[28866]=38027;
squeal_samples[28867]=39552;
squeal_samples[28868]=41020;
squeal_samples[28869]=42409;
squeal_samples[28870]=43744;
squeal_samples[28871]=45016;
squeal_samples[28872]=46232;
squeal_samples[28873]=47396;
squeal_samples[28874]=48500;
squeal_samples[28875]=49562;
squeal_samples[28876]=50570;
squeal_samples[28877]=51539;
squeal_samples[28878]=52458;
squeal_samples[28879]=53340;
squeal_samples[28880]=54186;
squeal_samples[28881]=52405;
squeal_samples[28882]=46718;
squeal_samples[28883]=41335;
squeal_samples[28884]=36311;
squeal_samples[28885]=31594;
squeal_samples[28886]=27186;
squeal_samples[28887]=23058;
squeal_samples[28888]=19205;
squeal_samples[28889]=15585;
squeal_samples[28890]=12206;
squeal_samples[28891]=9041;
squeal_samples[28892]=6079;
squeal_samples[28893]=4928;
squeal_samples[28894]=7739;
squeal_samples[28895]=10608;
squeal_samples[28896]=13354;
squeal_samples[28897]=15979;
squeal_samples[28898]=18490;
squeal_samples[28899]=20885;
squeal_samples[28900]=23177;
squeal_samples[28901]=25377;
squeal_samples[28902]=27464;
squeal_samples[28903]=29473;
squeal_samples[28904]=31379;
squeal_samples[28905]=33209;
squeal_samples[28906]=34952;
squeal_samples[28907]=36621;
squeal_samples[28908]=38213;
squeal_samples[28909]=39731;
squeal_samples[28910]=41185;
squeal_samples[28911]=42576;
squeal_samples[28912]=43897;
squeal_samples[28913]=45164;
squeal_samples[28914]=46368;
squeal_samples[28915]=47524;
squeal_samples[28916]=48627;
squeal_samples[28917]=49679;
squeal_samples[28918]=50686;
squeal_samples[28919]=51647;
squeal_samples[28920]=52560;
squeal_samples[28921]=53438;
squeal_samples[28922]=54279;
squeal_samples[28923]=51710;
squeal_samples[28924]=46014;
squeal_samples[28925]=40682;
squeal_samples[28926]=35686;
squeal_samples[28927]=31022;
squeal_samples[28928]=26642;
squeal_samples[28929]=22551;
squeal_samples[28930]=18728;
squeal_samples[28931]=15140;
squeal_samples[28932]=11790;
squeal_samples[28933]=8653;
squeal_samples[28934]=5713;
squeal_samples[28935]=5162;
squeal_samples[28936]=8096;
squeal_samples[28937]=10952;
squeal_samples[28938]=13677;
squeal_samples[28939]=16290;
squeal_samples[28940]=18790;
squeal_samples[28941]=21162;
squeal_samples[28942]=23449;
squeal_samples[28943]=25625;
squeal_samples[28944]=27714;
squeal_samples[28945]=29701;
squeal_samples[28946]=31605;
squeal_samples[28947]=33418;
squeal_samples[28948]=35159;
squeal_samples[28949]=36811;
squeal_samples[28950]=38396;
squeal_samples[28951]=39905;
squeal_samples[28952]=41353;
squeal_samples[28953]=42732;
squeal_samples[28954]=44044;
squeal_samples[28955]=45306;
squeal_samples[28956]=46505;
squeal_samples[28957]=47658;
squeal_samples[28958]=48749;
squeal_samples[28959]=49794;
squeal_samples[28960]=50793;
squeal_samples[28961]=51750;
squeal_samples[28962]=52663;
squeal_samples[28963]=53537;
squeal_samples[28964]=54317;
squeal_samples[28965]=50968;
squeal_samples[28966]=45323;
squeal_samples[28967]=40024;
squeal_samples[28968]=35083;
squeal_samples[28969]=30443;
squeal_samples[28970]=26103;
squeal_samples[28971]=22050;
squeal_samples[28972]=18251;
squeal_samples[28973]=14702;
squeal_samples[28974]=11373;
squeal_samples[28975]=8256;
squeal_samples[28976]=5355;
squeal_samples[28977]=5476;
squeal_samples[28978]=8455;
squeal_samples[28979]=11284;
squeal_samples[28980]=14000;
squeal_samples[28981]=16598;
squeal_samples[28982]=19082;
squeal_samples[28983]=21447;
squeal_samples[28984]=23716;
squeal_samples[28985]=25884;
squeal_samples[28986]=27953;
squeal_samples[28987]=29934;
squeal_samples[28988]=31822;
squeal_samples[28989]=33633;
squeal_samples[28990]=35358;
squeal_samples[28991]=36999;
squeal_samples[28992]=38578;
squeal_samples[28993]=40074;
squeal_samples[28994]=41520;
squeal_samples[28995]=42885;
squeal_samples[28996]=44199;
squeal_samples[28997]=45443;
squeal_samples[28998]=46640;
squeal_samples[28999]=47783;
squeal_samples[29000]=48871;
squeal_samples[29001]=49912;
squeal_samples[29002]=50907;
squeal_samples[29003]=51854;
squeal_samples[29004]=52761;
squeal_samples[29005]=53633;
squeal_samples[29006]=54247;
squeal_samples[29007]=50230;
squeal_samples[29008]=44625;
squeal_samples[29009]=39380;
squeal_samples[29010]=34474;
squeal_samples[29011]=29870;
squeal_samples[29012]=25574;
squeal_samples[29013]=21547;
squeal_samples[29014]=17786;
squeal_samples[29015]=14261;
squeal_samples[29016]=10964;
squeal_samples[29017]=7879;
squeal_samples[29018]=5033;
squeal_samples[29019]=5853;
squeal_samples[29020]=8795;
squeal_samples[29021]=11622;
squeal_samples[29022]=14315;
squeal_samples[29023]=16905;
squeal_samples[29024]=19366;
squeal_samples[29025]=21726;
squeal_samples[29026]=23981;
squeal_samples[29027]=26139;
squeal_samples[29028]=28191;
squeal_samples[29029]=30167;
squeal_samples[29030]=32039;
squeal_samples[29031]=33840;
squeal_samples[29032]=35551;
squeal_samples[29033]=37190;
squeal_samples[29034]=38761;
squeal_samples[29035]=40249;
squeal_samples[29036]=41682;
squeal_samples[29037]=43036;
squeal_samples[29038]=44346;
squeal_samples[29039]=45583;
squeal_samples[29040]=46775;
squeal_samples[29041]=47909;
squeal_samples[29042]=48994;
squeal_samples[29043]=50027;
squeal_samples[29044]=51015;
squeal_samples[29045]=51963;
squeal_samples[29046]=52862;
squeal_samples[29047]=53728;
squeal_samples[29048]=54072;
squeal_samples[29049]=49496;
squeal_samples[29050]=43940;
squeal_samples[29051]=38740;
squeal_samples[29052]=33868;
squeal_samples[29053]=29314;
squeal_samples[29054]=25044;
squeal_samples[29055]=21054;
squeal_samples[29056]=17319;
squeal_samples[29057]=13825;
squeal_samples[29058]=10553;
squeal_samples[29059]=7489;
squeal_samples[29060]=4815;
squeal_samples[29061]=6211;
squeal_samples[29062]=9150;
squeal_samples[29063]=11952;
squeal_samples[29064]=14640;
squeal_samples[29065]=17205;
squeal_samples[29066]=19662;
squeal_samples[29067]=22000;
squeal_samples[29068]=24244;
squeal_samples[29069]=26384;
squeal_samples[29070]=28436;
squeal_samples[29071]=30387;
squeal_samples[29072]=32263;
squeal_samples[29073]=34039;
squeal_samples[29074]=35757;
squeal_samples[29075]=37377;
squeal_samples[29076]=38941;
squeal_samples[29077]=40421;
squeal_samples[29078]=41844;
squeal_samples[29079]=43194;
squeal_samples[29080]=44497;
squeal_samples[29081]=45726;
squeal_samples[29082]=46908;
squeal_samples[29083]=48039;
squeal_samples[29084]=49114;
squeal_samples[29085]=50139;
squeal_samples[29086]=51126;
squeal_samples[29087]=52063;
squeal_samples[29088]=52962;
squeal_samples[29089]=53819;
squeal_samples[29090]=53790;
squeal_samples[29091]=48774;
squeal_samples[29092]=43259;
squeal_samples[29093]=38099;
squeal_samples[29094]=33271;
squeal_samples[29095]=28748;
squeal_samples[29096]=24519;
squeal_samples[29097]=20563;
squeal_samples[29098]=16864;
squeal_samples[29099]=13389;
squeal_samples[29100]=10151;
squeal_samples[29101]=7109;
squeal_samples[29102]=4683;
squeal_samples[29103]=6577;
squeal_samples[29104]=9495;
squeal_samples[29105]=12285;
squeal_samples[29106]=14952;
squeal_samples[29107]=17508;
squeal_samples[29108]=19945;
squeal_samples[29109]=22280;
squeal_samples[29110]=24507;
squeal_samples[29111]=26635;
squeal_samples[29112]=28673;
squeal_samples[29113]=30616;
squeal_samples[29114]=32479;
squeal_samples[29115]=34251;
squeal_samples[29116]=35951;
squeal_samples[29117]=37567;
squeal_samples[29118]=39118;
squeal_samples[29119]=40592;
squeal_samples[29120]=42004;
squeal_samples[29121]=43347;
squeal_samples[29122]=44644;
squeal_samples[29123]=45863;
squeal_samples[29124]=47042;
squeal_samples[29125]=48162;
squeal_samples[29126]=49233;
squeal_samples[29127]=50255;
squeal_samples[29128]=51232;
squeal_samples[29129]=52167;
squeal_samples[29130]=53060;
squeal_samples[29131]=53912;
squeal_samples[29132]=53404;
squeal_samples[29133]=48049;
squeal_samples[29134]=42589;
squeal_samples[29135]=37464;
squeal_samples[29136]=32683;
squeal_samples[29137]=28191;
squeal_samples[29138]=23997;
squeal_samples[29139]=20077;
squeal_samples[29140]=16398;
squeal_samples[29141]=12963;
squeal_samples[29142]=9746;
squeal_samples[29143]=6736;
squeal_samples[29144]=4642;
squeal_samples[29145]=6938;
squeal_samples[29146]=9840;
squeal_samples[29147]=12613;
squeal_samples[29148]=15266;
squeal_samples[29149]=17810;
squeal_samples[29150]=20234;
squeal_samples[29151]=22551;
squeal_samples[29152]=24766;
squeal_samples[29153]=26887;
squeal_samples[29154]=28907;
squeal_samples[29155]=30848;
squeal_samples[29156]=32692;
squeal_samples[29157]=34455;
squeal_samples[29158]=36143;
squeal_samples[29159]=37753;
squeal_samples[29160]=39290;
squeal_samples[29161]=40762;
squeal_samples[29162]=42163;
squeal_samples[29163]=43509;
squeal_samples[29164]=44783;
squeal_samples[29165]=46011;
squeal_samples[29166]=47172;
squeal_samples[29167]=48289;
squeal_samples[29168]=49353;
squeal_samples[29169]=50364;
squeal_samples[29170]=51345;
squeal_samples[29171]=52265;
squeal_samples[29172]=53162;
squeal_samples[29173]=53999;
squeal_samples[29174]=53494;
squeal_samples[29175]=48129;
squeal_samples[29176]=42662;
squeal_samples[29177]=37540;
squeal_samples[29178]=32740;
squeal_samples[29179]=28258;
squeal_samples[29180]=24050;
squeal_samples[29181]=20135;
squeal_samples[29182]=16445;
squeal_samples[29183]=13006;
squeal_samples[29184]=9785;
squeal_samples[29185]=6770;
squeal_samples[29186]=4679;
squeal_samples[29187]=6966;
squeal_samples[29188]=9871;
squeal_samples[29189]=12640;
squeal_samples[29190]=15296;
squeal_samples[29191]=17830;
squeal_samples[29192]=20257;
squeal_samples[29193]=22570;
squeal_samples[29194]=24783;
squeal_samples[29195]=26907;
squeal_samples[29196]=28925;
squeal_samples[29197]=30864;
squeal_samples[29198]=32705;
squeal_samples[29199]=34473;
squeal_samples[29200]=36158;
squeal_samples[29201]=37765;
squeal_samples[29202]=39300;
squeal_samples[29203]=40772;
squeal_samples[29204]=42168;
squeal_samples[29205]=43514;
squeal_samples[29206]=44789;
squeal_samples[29207]=46014;
squeal_samples[29208]=47180;
squeal_samples[29209]=48292;
squeal_samples[29210]=49357;
squeal_samples[29211]=50374;
squeal_samples[29212]=51342;
squeal_samples[29213]=52274;
squeal_samples[29214]=53154;
squeal_samples[29215]=54009;
squeal_samples[29216]=53491;
squeal_samples[29217]=48129;
squeal_samples[29218]=42664;
squeal_samples[29219]=37530;
squeal_samples[29220]=32739;
squeal_samples[29221]=28253;
squeal_samples[29222]=24048;
squeal_samples[29223]=20126;
squeal_samples[29224]=16442;
squeal_samples[29225]=12997;
squeal_samples[29226]=9788;
squeal_samples[29227]=6763;
squeal_samples[29228]=4672;
squeal_samples[29229]=6962;
squeal_samples[29230]=9863;
squeal_samples[29231]=12632;
squeal_samples[29232]=15289;
squeal_samples[29233]=17823;
squeal_samples[29234]=20254;
squeal_samples[29235]=22561;
squeal_samples[29236]=24781;
squeal_samples[29237]=26894;
squeal_samples[29238]=28920;
squeal_samples[29239]=30852;
squeal_samples[29240]=32694;
squeal_samples[29241]=34463;
squeal_samples[29242]=36145;
squeal_samples[29243]=37761;
squeal_samples[29244]=39294;
squeal_samples[29245]=40759;
squeal_samples[29246]=42165;
squeal_samples[29247]=43506;
squeal_samples[29248]=44779;
squeal_samples[29249]=46003;
squeal_samples[29250]=47168;
squeal_samples[29251]=48281;
squeal_samples[29252]=49347;
squeal_samples[29253]=50361;
squeal_samples[29254]=51334;
squeal_samples[29255]=52265;
squeal_samples[29256]=53144;
squeal_samples[29257]=54000;
squeal_samples[29258]=53476;
squeal_samples[29259]=48123;
squeal_samples[29260]=42647;
squeal_samples[29261]=37529;
squeal_samples[29262]=32732;
squeal_samples[29263]=28241;
squeal_samples[29264]=24040;
squeal_samples[29265]=20111;
squeal_samples[29266]=16433;
squeal_samples[29267]=12992;
squeal_samples[29268]=9774;
squeal_samples[29269]=6756;
squeal_samples[29270]=4657;
squeal_samples[29271]=6954;
squeal_samples[29272]=9849;
squeal_samples[29273]=12624;
squeal_samples[29274]=15275;
squeal_samples[29275]=17814;
squeal_samples[29276]=20240;
squeal_samples[29277]=22553;
squeal_samples[29278]=24767;
squeal_samples[29279]=26886;
squeal_samples[29280]=28906;
squeal_samples[29281]=30842;
squeal_samples[29282]=32684;
squeal_samples[29283]=34456;
squeal_samples[29284]=36134;
squeal_samples[29285]=37751;
squeal_samples[29286]=39281;
squeal_samples[29287]=40749;
squeal_samples[29288]=42154;
squeal_samples[29289]=43493;
squeal_samples[29290]=44772;
squeal_samples[29291]=45988;
squeal_samples[29292]=47159;
squeal_samples[29293]=48269;
squeal_samples[29294]=49335;
squeal_samples[29295]=50352;
squeal_samples[29296]=51321;
squeal_samples[29297]=52255;
squeal_samples[29298]=53134;
squeal_samples[29299]=53985;
squeal_samples[29300]=53470;
squeal_samples[29301]=48107;
squeal_samples[29302]=42640;
squeal_samples[29303]=37515;
squeal_samples[29304]=32723;
squeal_samples[29305]=28228;
squeal_samples[29306]=24029;
squeal_samples[29307]=20102;
squeal_samples[29308]=16424;
squeal_samples[29309]=12985;
squeal_samples[29310]=9759;
squeal_samples[29311]=6747;
squeal_samples[29312]=4646;
squeal_samples[29313]=6941;
squeal_samples[29314]=9841;
squeal_samples[29315]=12609;
squeal_samples[29316]=15267;
squeal_samples[29317]=17803;
squeal_samples[29318]=20227;
squeal_samples[29319]=22544;
squeal_samples[29320]=24754;
squeal_samples[29321]=26876;
squeal_samples[29322]=28894;
squeal_samples[29323]=30833;
squeal_samples[29324]=32676;
squeal_samples[29325]=34446;
squeal_samples[29326]=36123;
squeal_samples[29327]=37739;
squeal_samples[29328]=39270;
squeal_samples[29329]=40739;
squeal_samples[29330]=42143;
squeal_samples[29331]=43481;
squeal_samples[29332]=44761;
squeal_samples[29333]=45977;
squeal_samples[29334]=47148;
squeal_samples[29335]=48258;
squeal_samples[29336]=49325;
squeal_samples[29337]=50338;
squeal_samples[29338]=51314;
squeal_samples[29339]=52240;
squeal_samples[29340]=53125;
squeal_samples[29341]=53974;
squeal_samples[29342]=53457;
squeal_samples[29343]=48099;
squeal_samples[29344]=42626;
squeal_samples[29345]=37505;
squeal_samples[29346]=32711;
squeal_samples[29347]=28219;
squeal_samples[29348]=24015;
squeal_samples[29349]=20094;
squeal_samples[29350]=16411;
squeal_samples[29351]=12973;
squeal_samples[29352]=9751;
squeal_samples[29353]=6733;
squeal_samples[29354]=4636;
squeal_samples[29355]=6932;
squeal_samples[29356]=9826;
squeal_samples[29357]=12602;
squeal_samples[29358]=15253;
squeal_samples[29359]=17792;
squeal_samples[29360]=20219;
squeal_samples[29361]=22529;
squeal_samples[29362]=24747;
squeal_samples[29363]=26860;
squeal_samples[29364]=28887;
squeal_samples[29365]=30819;
squeal_samples[29366]=32668;
squeal_samples[29367]=34432;
squeal_samples[29368]=36115;
squeal_samples[29369]=37723;
squeal_samples[29370]=39266;
squeal_samples[29371]=40721;
squeal_samples[29372]=42137;
squeal_samples[29373]=43468;
squeal_samples[29374]=44749;
squeal_samples[29375]=45968;
squeal_samples[29376]=47135;
squeal_samples[29377]=48249;
squeal_samples[29378]=49312;
squeal_samples[29379]=50329;
squeal_samples[29380]=51301;
squeal_samples[29381]=52230;
squeal_samples[29382]=53114;
squeal_samples[29383]=53961;
squeal_samples[29384]=53450;
squeal_samples[29385]=48083;
squeal_samples[29386]=42619;
squeal_samples[29387]=37492;
squeal_samples[29388]=32701;
squeal_samples[29389]=28207;
squeal_samples[29390]=24006;
squeal_samples[29391]=20079;
squeal_samples[29392]=16404;
squeal_samples[29393]=12961;
squeal_samples[29394]=9738;
squeal_samples[29395]=6726;
squeal_samples[29396]=4620;
squeal_samples[29397]=6925;
squeal_samples[29398]=9813;
squeal_samples[29399]=12592;
squeal_samples[29400]=15240;
squeal_samples[29401]=17784;
squeal_samples[29402]=20203;
squeal_samples[29403]=22525;
squeal_samples[29404]=24729;
squeal_samples[29405]=26855;
squeal_samples[29406]=28871;
squeal_samples[29407]=30811;
squeal_samples[29408]=32655;
squeal_samples[29409]=34423;
squeal_samples[29410]=36102;
squeal_samples[29411]=37715;
squeal_samples[29412]=39250;
squeal_samples[29413]=40715;
squeal_samples[29414]=42121;
squeal_samples[29415]=43462;
squeal_samples[29416]=44734;
squeal_samples[29417]=45960;
squeal_samples[29418]=47121;
squeal_samples[29419]=48241;
squeal_samples[29420]=49298;
squeal_samples[29421]=50320;
squeal_samples[29422]=51288;
squeal_samples[29423]=52222;
squeal_samples[29424]=53100;
squeal_samples[29425]=53953;
squeal_samples[29426]=53435;
squeal_samples[29427]=48076;
squeal_samples[29428]=42605;
squeal_samples[29429]=37483;
squeal_samples[29430]=32688;
squeal_samples[29431]=28197;
squeal_samples[29432]=23995;
squeal_samples[29433]=20068;
squeal_samples[29434]=16393;
squeal_samples[29435]=12949;
squeal_samples[29436]=9729;
squeal_samples[29437]=6711;
squeal_samples[29438]=4615;
squeal_samples[29439]=6906;
squeal_samples[29440]=9810;
squeal_samples[29441]=12574;
squeal_samples[29442]=15236;
squeal_samples[29443]=17767;
squeal_samples[29444]=20197;
squeal_samples[29445]=22508;
squeal_samples[29446]=24724;
squeal_samples[29447]=26839;
squeal_samples[29448]=28864;
squeal_samples[29449]=30798;
squeal_samples[29450]=32643;
squeal_samples[29451]=34415;
squeal_samples[29452]=36087;
squeal_samples[29453]=37708;
squeal_samples[29454]=39236;
squeal_samples[29455]=40706;
squeal_samples[29456]=42109;
squeal_samples[29457]=43450;
squeal_samples[29458]=44725;
squeal_samples[29459]=45947;
squeal_samples[29460]=47112;
squeal_samples[29461]=48227;
squeal_samples[29462]=49291;
squeal_samples[29463]=50305;
squeal_samples[29464]=51279;
squeal_samples[29465]=52210;
squeal_samples[29466]=53089;
squeal_samples[29467]=53943;
squeal_samples[29468]=53423;
squeal_samples[29469]=48065;
squeal_samples[29470]=42594;
squeal_samples[29471]=37472;
squeal_samples[29472]=32677;
squeal_samples[29473]=28186;
squeal_samples[29474]=23984;
squeal_samples[29475]=20056;
squeal_samples[29476]=16383;
squeal_samples[29477]=12937;
squeal_samples[29478]=9719;
squeal_samples[29479]=6699;
squeal_samples[29480]=4604;
squeal_samples[29481]=6896;
squeal_samples[29482]=9798;
squeal_samples[29483]=12564;
squeal_samples[29484]=15222;
squeal_samples[29485]=17759;
squeal_samples[29486]=20185;
squeal_samples[29487]=22497;
squeal_samples[29488]=24713;
squeal_samples[29489]=26827;
squeal_samples[29490]=28855;
squeal_samples[29491]=30784;
squeal_samples[29492]=32635;
squeal_samples[29493]=34401;
squeal_samples[29494]=36079;
squeal_samples[29495]=37694;
squeal_samples[29496]=39227;
squeal_samples[29497]=40693;
squeal_samples[29498]=42099;
squeal_samples[29499]=43440;
squeal_samples[29500]=44711;
squeal_samples[29501]=45938;
squeal_samples[29502]=47100;
squeal_samples[29503]=48216;
squeal_samples[29504]=49280;
squeal_samples[29505]=50294;
squeal_samples[29506]=51267;
squeal_samples[29507]=52199;
squeal_samples[29508]=53077;
squeal_samples[29509]=53932;
squeal_samples[29510]=53889;
squeal_samples[29511]=48860;
squeal_samples[29512]=43330;
squeal_samples[29513]=38163;
squeal_samples[29514]=33322;
squeal_samples[29515]=28789;
squeal_samples[29516]=24549;
squeal_samples[29517]=20577;
squeal_samples[29518]=16871;
squeal_samples[29519]=13398;
squeal_samples[29520]=10148;
squeal_samples[29521]=7102;
squeal_samples[29522]=4668;
squeal_samples[29523]=6554;
squeal_samples[29524]=9469;
squeal_samples[29525]=12256;
squeal_samples[29526]=14923;
squeal_samples[29527]=17470;
squeal_samples[29528]=19908;
squeal_samples[29529]=22237;
squeal_samples[29530]=24461;
squeal_samples[29531]=26590;
squeal_samples[29532]=28625;
squeal_samples[29533]=30568;
squeal_samples[29534]=32425;
squeal_samples[29535]=34189;
squeal_samples[29536]=35889;
squeal_samples[29537]=37499;
squeal_samples[29538]=39052;
squeal_samples[29539]=40523;
squeal_samples[29540]=41936;
squeal_samples[29541]=43280;
squeal_samples[29542]=44569;
squeal_samples[29543]=45792;
squeal_samples[29544]=46968;
squeal_samples[29545]=48083;
squeal_samples[29546]=49155;
squeal_samples[29547]=50175;
squeal_samples[29548]=51153;
squeal_samples[29549]=52084;
squeal_samples[29550]=52974;
squeal_samples[29551]=53828;
squeal_samples[29552]=54159;
squeal_samples[29553]=49578;
squeal_samples[29554]=43997;
squeal_samples[29555]=38790;
squeal_samples[29556]=33905;
squeal_samples[29557]=29341;
squeal_samples[29558]=25060;
squeal_samples[29559]=21064;
squeal_samples[29560]=17318;
squeal_samples[29561]=13814;
squeal_samples[29562]=10536;
squeal_samples[29563]=7469;
squeal_samples[29564]=4779;
squeal_samples[29565]=6181;
squeal_samples[29566]=9104;
squeal_samples[29567]=11908;
squeal_samples[29568]=14593;
squeal_samples[29569]=17153;
squeal_samples[29570]=19605;
squeal_samples[29571]=21943;
squeal_samples[29572]=24181;
squeal_samples[29573]=26321;
squeal_samples[29574]=28368;
squeal_samples[29575]=30314;
squeal_samples[29576]=32188;
squeal_samples[29577]=33968;
squeal_samples[29578]=35675;
squeal_samples[29579]=37295;
squeal_samples[29580]=38855;
squeal_samples[29581]=40332;
squeal_samples[29582]=41753;
squeal_samples[29583]=43106;
squeal_samples[29584]=44400;
squeal_samples[29585]=45636;
squeal_samples[29586]=46814;
squeal_samples[29587]=47938;
squeal_samples[29588]=49012;
squeal_samples[29589]=50040;
squeal_samples[29590]=51023;
squeal_samples[29591]=51957;
squeal_samples[29592]=52857;
squeal_samples[29593]=53709;
squeal_samples[29594]=54322;
squeal_samples[29595]=50284;
squeal_samples[29596]=44671;
squeal_samples[29597]=39408;
squeal_samples[29598]=34492;
squeal_samples[29599]=29884;
squeal_samples[29600]=25570;
squeal_samples[29601]=21531;
squeal_samples[29602]=17769;
squeal_samples[29603]=14227;
squeal_samples[29604]=10926;
squeal_samples[29605]=7828;
squeal_samples[29606]=4985;
squeal_samples[29607]=5790;
squeal_samples[29608]=8738;
squeal_samples[29609]=11554;
squeal_samples[29610]=14249;
squeal_samples[29611]=16830;
squeal_samples[29612]=19293;
squeal_samples[29613]=21645;
squeal_samples[29614]=23898;
squeal_samples[29615]=26046;
squeal_samples[29616]=28105;
squeal_samples[29617]=30066;
squeal_samples[29618]=31948;
squeal_samples[29619]=33741;
squeal_samples[29620]=35451;
squeal_samples[29621]=37090;
squeal_samples[29622]=38652;
squeal_samples[29623]=40145;
squeal_samples[29624]=41566;
squeal_samples[29625]=42929;
squeal_samples[29626]=44229;
squeal_samples[29627]=45476;
squeal_samples[29628]=46653;
squeal_samples[29629]=47794;
squeal_samples[29630]=48870;
squeal_samples[29631]=49905;
squeal_samples[29632]=50891;
squeal_samples[29633]=51833;
squeal_samples[29634]=52735;
squeal_samples[29635]=53598;
squeal_samples[29636]=54365;
squeal_samples[29637]=51008;
squeal_samples[29638]=45337;
squeal_samples[29639]=40046;
squeal_samples[29640]=35072;
squeal_samples[29641]=30435;
squeal_samples[29642]=26086;
squeal_samples[29643]=22007;
squeal_samples[29644]=18216;
squeal_samples[29645]=14644;
squeal_samples[29646]=11318;
squeal_samples[29647]=8192;
squeal_samples[29648]=5278;
squeal_samples[29649]=5399;
squeal_samples[29650]=8366;
squeal_samples[29651]=11198;
squeal_samples[29652]=13905;
squeal_samples[29653]=16505;
squeal_samples[29654]=18978;
squeal_samples[29655]=21345;
squeal_samples[29656]=23612;
squeal_samples[29657]=25773;
squeal_samples[29658]=27845;
squeal_samples[29659]=29817;
squeal_samples[29660]=31708;
squeal_samples[29661]=33508;
squeal_samples[29662]=35235;
squeal_samples[29663]=36877;
squeal_samples[29664]=38447;
squeal_samples[29665]=39949;
squeal_samples[29666]=41381;
squeal_samples[29667]=42756;
squeal_samples[29668]=44061;
squeal_samples[29669]=45311;
squeal_samples[29670]=46499;
squeal_samples[29671]=47639;
squeal_samples[29672]=48730;
squeal_samples[29673]=49768;
squeal_samples[29674]=50762;
squeal_samples[29675]=51706;
squeal_samples[29676]=52618;
squeal_samples[29677]=53480;
squeal_samples[29678]=54309;
squeal_samples[29679]=51725;
squeal_samples[29680]=46018;
squeal_samples[29681]=40668;
squeal_samples[29682]=35670;
squeal_samples[29683]=30981;
squeal_samples[29684]=26601;
squeal_samples[29685]=22494;
squeal_samples[29686]=18662;
squeal_samples[29687]=15072;
squeal_samples[29688]=11709;
squeal_samples[29689]=8567;
squeal_samples[29690]=5616;
squeal_samples[29691]=5061;
squeal_samples[29692]=7988;
squeal_samples[29693]=10840;
squeal_samples[29694]=13563;
squeal_samples[29695]=16173;
squeal_samples[29696]=18664;
squeal_samples[29697]=21041;
squeal_samples[29698]=23323;
squeal_samples[29699]=25498;
squeal_samples[29700]=27578;
squeal_samples[29701]=29562;
squeal_samples[29702]=31464;
squeal_samples[29703]=33273;
squeal_samples[29704]=35014;
squeal_samples[29705]=36665;
squeal_samples[29706]=38246;
squeal_samples[29707]=39753;
squeal_samples[29708]=41198;
squeal_samples[29709]=42575;
squeal_samples[29710]=43889;
squeal_samples[29711]=45147;
squeal_samples[29712]=46348;
squeal_samples[29713]=47491;
squeal_samples[29714]=48585;
squeal_samples[29715]=49626;
squeal_samples[29716]=50625;
squeal_samples[29717]=51584;
squeal_samples[29718]=52489;
squeal_samples[29719]=53364;
squeal_samples[29720]=54195;
squeal_samples[29721]=52409;
squeal_samples[29722]=46699;
squeal_samples[29723]=41312;
squeal_samples[29724]=36265;
squeal_samples[29725]=31541;
squeal_samples[29726]=27121;
squeal_samples[29727]=22984;
squeal_samples[29728]=19117;
squeal_samples[29729]=15496;
squeal_samples[29730]=12106;
squeal_samples[29731]=8934;
squeal_samples[29732]=5967;
squeal_samples[29733]=4802;
squeal_samples[29734]=7616;
squeal_samples[29735]=10478;
squeal_samples[29736]=13224;
squeal_samples[29737]=15840;
squeal_samples[29738]=18349;
squeal_samples[29739]=20738;
squeal_samples[29740]=23028;
squeal_samples[29741]=25223;
squeal_samples[29742]=27310;
squeal_samples[29743]=29309;
squeal_samples[29744]=31219;
squeal_samples[29745]=33040;
squeal_samples[29746]=34790;
squeal_samples[29747]=36450;
squeal_samples[29748]=38037;
squeal_samples[29749]=39562;
squeal_samples[29750]=41003;
squeal_samples[29751]=42400;
squeal_samples[29752]=43712;
squeal_samples[29753]=44981;
squeal_samples[29754]=46183;
squeal_samples[29755]=47342;
squeal_samples[29756]=48435;
squeal_samples[29757]=49492;
squeal_samples[29758]=50495;
squeal_samples[29759]=51451;
squeal_samples[29760]=52374;
squeal_samples[29761]=53243;
squeal_samples[29762]=54087;
squeal_samples[29763]=52974;
squeal_samples[29764]=47393;
squeal_samples[29765]=41951;
squeal_samples[29766]=36868;
squeal_samples[29767]=32106;
squeal_samples[29768]=27648;
squeal_samples[29769]=23477;
squeal_samples[29770]=19581;
squeal_samples[29771]=15921;
squeal_samples[29772]=12507;
squeal_samples[29773]=9305;
squeal_samples[29774]=6318;
squeal_samples[29775]=4637;
squeal_samples[29776]=7235;
squeal_samples[29777]=10117;
squeal_samples[29778]=12872;
squeal_samples[29779]=15512;
squeal_samples[29780]=18027;
squeal_samples[29781]=20439;
squeal_samples[29782]=22744;
squeal_samples[29783]=24936;
squeal_samples[29784]=27048;
squeal_samples[29785]=29050;
squeal_samples[29786]=30977;
squeal_samples[29787]=32807;
squeal_samples[29788]=34562;
squeal_samples[29789]=36237;
squeal_samples[29790]=37833;
squeal_samples[29791]=39363;
squeal_samples[29792]=40823;
squeal_samples[29793]=42211;
squeal_samples[29794]=43547;
squeal_samples[29795]=44817;
squeal_samples[29796]=46026;
squeal_samples[29797]=47189;
squeal_samples[29798]=48295;
squeal_samples[29799]=49350;
squeal_samples[29800]=50359;
squeal_samples[29801]=51327;
squeal_samples[29802]=52247;
squeal_samples[29803]=53126;
squeal_samples[29804]=53970;
squeal_samples[29805]=53447;
squeal_samples[29806]=48084;
squeal_samples[29807]=42600;
squeal_samples[29808]=37475;
squeal_samples[29809]=32668;
squeal_samples[29810]=28181;
squeal_samples[29811]=23972;
squeal_samples[29812]=20039;
squeal_samples[29813]=16361;
squeal_samples[29814]=12908;
squeal_samples[29815]=9687;
squeal_samples[29816]=6664;
squeal_samples[29817]=4566;
squeal_samples[29818]=6858;
squeal_samples[29819]=9751;
squeal_samples[29820]=12529;
squeal_samples[29821]=15175;
squeal_samples[29822]=17711;
squeal_samples[29823]=20133;
squeal_samples[29824]=22449;
squeal_samples[29825]=24663;
squeal_samples[29826]=26772;
squeal_samples[29827]=28800;
squeal_samples[29828]=30728;
squeal_samples[29829]=32577;
squeal_samples[29830]=34337;
squeal_samples[29831]=36021;
squeal_samples[29832]=37627;
squeal_samples[29833]=39161;
squeal_samples[29834]=40634;
squeal_samples[29835]=42032;
squeal_samples[29836]=43372;
squeal_samples[29837]=44650;
squeal_samples[29838]=45867;
squeal_samples[29839]=47038;
squeal_samples[29840]=48148;
squeal_samples[29841]=49207;
squeal_samples[29842]=50225;
squeal_samples[29843]=51194;
squeal_samples[29844]=52123;
squeal_samples[29845]=53005;
squeal_samples[29846]=53854;
squeal_samples[29847]=54182;
squeal_samples[29848]=49591;
squeal_samples[29849]=44016;
squeal_samples[29850]=38797;
squeal_samples[29851]=33908;
squeal_samples[29852]=29336;
squeal_samples[29853]=25053;
squeal_samples[29854]=21043;
squeal_samples[29855]=17306;
squeal_samples[29856]=13794;
squeal_samples[29857]=10510;
squeal_samples[29858]=7439;
squeal_samples[29859]=4748;
squeal_samples[29860]=6146;
squeal_samples[29861]=9073;
squeal_samples[29862]=11868;
squeal_samples[29863]=14550;
squeal_samples[29864]=17108;
squeal_samples[29865]=19562;
squeal_samples[29866]=21899;
squeal_samples[29867]=24135;
squeal_samples[29868]=26275;
squeal_samples[29869]=28320;
squeal_samples[29870]=30268;
squeal_samples[29871]=32137;
squeal_samples[29872]=33913;
squeal_samples[29873]=35621;
squeal_samples[29874]=37245;
squeal_samples[29875]=38800;
squeal_samples[29876]=40278;
squeal_samples[29877]=41698;
squeal_samples[29878]=43046;
squeal_samples[29879]=44339;
squeal_samples[29880]=45576;
squeal_samples[29881]=46754;
squeal_samples[29882]=47877;
squeal_samples[29883]=48954;
squeal_samples[29884]=49976;
squeal_samples[29885]=50960;
squeal_samples[29886]=51894;
squeal_samples[29887]=52793;
squeal_samples[29888]=53642;
squeal_samples[29889]=54417;
squeal_samples[29890]=51042;
squeal_samples[29891]=45373;
squeal_samples[29892]=40068;
squeal_samples[29893]=35098;
squeal_samples[29894]=30443;
squeal_samples[29895]=26096;
squeal_samples[29896]=22015;
squeal_samples[29897]=18211;
squeal_samples[29898]=14643;
squeal_samples[29899]=11307;
squeal_samples[29900]=8186;
squeal_samples[29901]=5256;
squeal_samples[29902]=5388;
squeal_samples[29903]=8339;
squeal_samples[29904]=11179;
squeal_samples[29905]=13881;
squeal_samples[29906]=16479;
squeal_samples[29907]=18949;
squeal_samples[29908]=21314;
squeal_samples[29909]=23577;
squeal_samples[29910]=25742;
squeal_samples[29911]=27811;
squeal_samples[29912]=29784;
squeal_samples[29913]=31670;
squeal_samples[29914]=33469;
squeal_samples[29915]=35196;
squeal_samples[29916]=36841;
squeal_samples[29917]=38405;
squeal_samples[29918]=39908;
squeal_samples[29919]=41336;
squeal_samples[29920]=42712;
squeal_samples[29921]=44012;
squeal_samples[29922]=45262;
squeal_samples[29923]=46454;
squeal_samples[29924]=47591;
squeal_samples[29925]=48680;
squeal_samples[29926]=49719;
squeal_samples[29927]=50706;
squeal_samples[29928]=51659;
squeal_samples[29929]=52560;
squeal_samples[29930]=53428;
squeal_samples[29931]=54254;
squeal_samples[29932]=52459;
squeal_samples[29933]=46745;
squeal_samples[29934]=41352;
squeal_samples[29935]=36296;
squeal_samples[29936]=31568;
squeal_samples[29937]=27143;
squeal_samples[29938]=22999;
squeal_samples[29939]=19134;
squeal_samples[29940]=15505;
squeal_samples[29941]=12113;
squeal_samples[29942]=8932;
squeal_samples[29943]=5962;
squeal_samples[29944]=4797;
squeal_samples[29945]=7608;
squeal_samples[29946]=10470;
squeal_samples[29947]=13204;
squeal_samples[29948]=15831;
squeal_samples[29949]=18331;
squeal_samples[29950]=20722;
squeal_samples[29951]=23012;
squeal_samples[29952]=25201;
squeal_samples[29953]=27287;
squeal_samples[29954]=29288;
squeal_samples[29955]=31195;
squeal_samples[29956]=33021;
squeal_samples[29957]=34761;
squeal_samples[29958]=36423;
squeal_samples[29959]=38010;
squeal_samples[29960]=39533;
squeal_samples[29961]=40977;
squeal_samples[29962]=42366;
squeal_samples[29963]=43681;
squeal_samples[29964]=44947;
squeal_samples[29965]=46150;
squeal_samples[29966]=47303;
squeal_samples[29967]=48402;
squeal_samples[29968]=49456;
squeal_samples[29969]=50452;
squeal_samples[29970]=51419;
squeal_samples[29971]=52322;
squeal_samples[29972]=53206;
squeal_samples[29973]=54043;
squeal_samples[29974]=53514;
squeal_samples[29975]=48142;
squeal_samples[29976]=42650;
squeal_samples[29977]=37522;
squeal_samples[29978]=32712;
squeal_samples[29979]=28212;
squeal_samples[29980]=24006;
squeal_samples[29981]=20065;
squeal_samples[29982]=16377;
squeal_samples[29983]=12926;
squeal_samples[29984]=9697;
squeal_samples[29985]=6682;
squeal_samples[29986]=4571;
squeal_samples[29987]=6862;
squeal_samples[29988]=9753;
squeal_samples[29989]=12530;
squeal_samples[29990]=15169;
squeal_samples[29991]=17711;
squeal_samples[29992]=20127;
squeal_samples[29993]=22439;
squeal_samples[29994]=24650;
squeal_samples[29995]=26769;
squeal_samples[29996]=28787;
squeal_samples[29997]=30712;
squeal_samples[29998]=32560;
squeal_samples[29999]=34321;
squeal_samples[30000]=36005;
squeal_samples[30001]=37610;
squeal_samples[30002]=39145;
squeal_samples[30003]=40611;
squeal_samples[30004]=42010;
squeal_samples[30005]=43347;
squeal_samples[30006]=44624;
squeal_samples[30007]=45845;
squeal_samples[30008]=47005;
squeal_samples[30009]=48126;
squeal_samples[30010]=49176;
squeal_samples[30011]=50199;
squeal_samples[30012]=51167;
squeal_samples[30013]=52095;
squeal_samples[30014]=52979;
squeal_samples[30015]=53826;
squeal_samples[30016]=54154;
squeal_samples[30017]=49559;
squeal_samples[30018]=43984;
squeal_samples[30019]=38763;
squeal_samples[30020]=33875;
squeal_samples[30021]=29300;
squeal_samples[30022]=25016;
squeal_samples[30023]=21016;
squeal_samples[30024]=17264;
squeal_samples[30025]=13755;
squeal_samples[30026]=10475;
squeal_samples[30027]=7397;
squeal_samples[30028]=4714;
squeal_samples[30029]=6105;
squeal_samples[30030]=9036;
squeal_samples[30031]=11830;
squeal_samples[30032]=14510;
squeal_samples[30033]=17073;
squeal_samples[30034]=19522;
squeal_samples[30035]=21860;
squeal_samples[30036]=24100;
squeal_samples[30037]=26233;
squeal_samples[30038]=28280;
squeal_samples[30039]=30228;
squeal_samples[30040]=32099;
squeal_samples[30041]=33876;
squeal_samples[30042]=35581;
squeal_samples[30043]=37203;
squeal_samples[30044]=38756;
squeal_samples[30045]=40240;
squeal_samples[30046]=41659;
squeal_samples[30047]=43009;
squeal_samples[30048]=44299;
squeal_samples[30049]=45536;
squeal_samples[30050]=46706;
squeal_samples[30051]=47838;
squeal_samples[30052]=48906;
squeal_samples[30053]=49936;
squeal_samples[30054]=50920;
squeal_samples[30055]=51851;
squeal_samples[30056]=52756;
squeal_samples[30057]=53602;
squeal_samples[30058]=54376;
squeal_samples[30059]=51001;
squeal_samples[30060]=45333;
squeal_samples[30061]=40021;
squeal_samples[30062]=35056;
squeal_samples[30063]=30405;
squeal_samples[30064]=26052;
squeal_samples[30065]=21977;
squeal_samples[30066]=18168;
squeal_samples[30067]=14599;
squeal_samples[30068]=11264;
squeal_samples[30069]=8141;
squeal_samples[30070]=5215;
squeal_samples[30071]=5342;
squeal_samples[30072]=8299;
squeal_samples[30073]=11131;
squeal_samples[30074]=13842;
squeal_samples[30075]=16432;
squeal_samples[30076]=18909;
squeal_samples[30077]=21273;
squeal_samples[30078]=23534;
squeal_samples[30079]=25699;
squeal_samples[30080]=27767;
squeal_samples[30081]=29741;
squeal_samples[30082]=31626;
squeal_samples[30083]=33426;
squeal_samples[30084]=35153;
squeal_samples[30085]=36795;
squeal_samples[30086]=38365;
squeal_samples[30087]=39861;
squeal_samples[30088]=41296;
squeal_samples[30089]=42666;
squeal_samples[30090]=43970;
squeal_samples[30091]=45216;
squeal_samples[30092]=46414;
squeal_samples[30093]=47550;
squeal_samples[30094]=48638;
squeal_samples[30095]=49675;
squeal_samples[30096]=50662;
squeal_samples[30097]=51616;
squeal_samples[30098]=52517;
squeal_samples[30099]=53383;
squeal_samples[30100]=54212;
squeal_samples[30101]=52415;
squeal_samples[30102]=46701;
squeal_samples[30103]=41309;
squeal_samples[30104]=36253;
squeal_samples[30105]=31523;
squeal_samples[30106]=27102;
squeal_samples[30107]=22958;
squeal_samples[30108]=19092;
squeal_samples[30109]=15462;
squeal_samples[30110]=12068;
squeal_samples[30111]=8890;
squeal_samples[30112]=5917;
squeal_samples[30113]=4754;
squeal_samples[30114]=7566;
squeal_samples[30115]=10424;
squeal_samples[30116]=13168;
squeal_samples[30117]=15785;
squeal_samples[30118]=18290;
squeal_samples[30119]=20677;
squeal_samples[30120]=22970;
squeal_samples[30121]=25154;
squeal_samples[30122]=27247;
squeal_samples[30123]=29242;
squeal_samples[30124]=31153;
squeal_samples[30125]=32976;
squeal_samples[30126]=34717;
squeal_samples[30127]=36380;
squeal_samples[30128]=37966;
squeal_samples[30129]=39491;
squeal_samples[30130]=40931;
squeal_samples[30131]=42324;
squeal_samples[30132]=43635;
squeal_samples[30133]=44905;
squeal_samples[30134]=46108;
squeal_samples[30135]=47256;
squeal_samples[30136]=48364;
squeal_samples[30137]=49403;
squeal_samples[30138]=50419;
squeal_samples[30139]=51366;
squeal_samples[30140]=52285;
squeal_samples[30141]=53160;
squeal_samples[30142]=53998;
squeal_samples[30143]=53474;
squeal_samples[30144]=48094;
squeal_samples[30145]=42610;
squeal_samples[30146]=37475;
squeal_samples[30147]=32671;
squeal_samples[30148]=28169;
squeal_samples[30149]=23959;
squeal_samples[30150]=20025;
squeal_samples[30151]=16330;
squeal_samples[30152]=12883;
squeal_samples[30153]=9657;
squeal_samples[30154]=6635;
squeal_samples[30155]=4528;
squeal_samples[30156]=6819;
squeal_samples[30157]=9708;
squeal_samples[30158]=12487;
squeal_samples[30159]=15126;
squeal_samples[30160]=17666;
squeal_samples[30161]=20085;
squeal_samples[30162]=22394;
squeal_samples[30163]=24607;
squeal_samples[30164]=26724;
squeal_samples[30165]=28745;
squeal_samples[30166]=30667;
squeal_samples[30167]=32517;
squeal_samples[30168]=34278;
squeal_samples[30169]=35960;
squeal_samples[30170]=37567;
squeal_samples[30171]=39100;
squeal_samples[30172]=40569;
squeal_samples[30173]=41965;
squeal_samples[30174]=43304;
squeal_samples[30175]=44580;
squeal_samples[30176]=45800;
squeal_samples[30177]=46964;
squeal_samples[30178]=48077;
squeal_samples[30179]=49138;
squeal_samples[30180]=50151;
squeal_samples[30181]=51126;
squeal_samples[30182]=52049;
squeal_samples[30183]=52934;
squeal_samples[30184]=53783;
squeal_samples[30185]=54376;
squeal_samples[30186]=50330;
squeal_samples[30187]=44701;
squeal_samples[30188]=39429;
squeal_samples[30189]=34501;
squeal_samples[30190]=29885;
squeal_samples[30191]=25560;
squeal_samples[30192]=21519;
squeal_samples[30193]=17736;
squeal_samples[30194]=14191;
squeal_samples[30195]=10880;
squeal_samples[30196]=7779;
squeal_samples[30197]=4924;
squeal_samples[30198]=5730;
squeal_samples[30199]=8671;
squeal_samples[30200]=11482;
squeal_samples[30201]=14179;
squeal_samples[30202]=16751;
squeal_samples[30203]=19213;
squeal_samples[30204]=21560;
squeal_samples[30205]=23812;
squeal_samples[30206]=25958;
squeal_samples[30207]=28010;
squeal_samples[30208]=29976;
squeal_samples[30209]=31845;
squeal_samples[30210]=33641;
squeal_samples[30211]=35349;
squeal_samples[30212]=36989;
squeal_samples[30213]=38539;
squeal_samples[30214]=40038;
squeal_samples[30215]=41455;
squeal_samples[30216]=42819;
squeal_samples[30217]=44117;
squeal_samples[30218]=45350;
squeal_samples[30219]=46544;
squeal_samples[30220]=47668;
squeal_samples[30221]=48753;
squeal_samples[30222]=49782;
squeal_samples[30223]=50765;
squeal_samples[30224]=51708;
squeal_samples[30225]=52607;
squeal_samples[30226]=53471;
squeal_samples[30227]=54289;
squeal_samples[30228]=52486;
squeal_samples[30229]=46770;
squeal_samples[30230]=41365;
squeal_samples[30231]=36307;
squeal_samples[30232]=31574;
squeal_samples[30233]=27142;
squeal_samples[30234]=22997;
squeal_samples[30235]=19125;
squeal_samples[30236]=15486;
squeal_samples[30237]=12091;
squeal_samples[30238]=8911;
squeal_samples[30239]=5938;
squeal_samples[30240]=4770;
squeal_samples[30241]=7576;
squeal_samples[30242]=10434;
squeal_samples[30243]=13174;
squeal_samples[30244]=15789;
squeal_samples[30245]=18295;
squeal_samples[30246]=20682;
squeal_samples[30247]=22969;
squeal_samples[30248]=25156;
squeal_samples[30249]=27242;
squeal_samples[30250]=29246;
squeal_samples[30251]=31144;
squeal_samples[30252]=32972;
squeal_samples[30253]=34711;
squeal_samples[30254]=36372;
squeal_samples[30255]=37957;
squeal_samples[30256]=39476;
squeal_samples[30257]=40926;
squeal_samples[30258]=42306;
squeal_samples[30259]=43628;
squeal_samples[30260]=44886;
squeal_samples[30261]=46090;
squeal_samples[30262]=47242;
squeal_samples[30263]=48343;
squeal_samples[30264]=49392;
squeal_samples[30265]=50390;
squeal_samples[30266]=51355;
squeal_samples[30267]=52263;
squeal_samples[30268]=53145;
squeal_samples[30269]=53976;
squeal_samples[30270]=53926;
squeal_samples[30271]=48880;
squeal_samples[30272]=43339;
squeal_samples[30273]=38157;
squeal_samples[30274]=33303;
squeal_samples[30275]=28760;
squeal_samples[30276]=24508;
squeal_samples[30277]=20534;
squeal_samples[30278]=16813;
squeal_samples[30279]=13329;
squeal_samples[30280]=10067;
squeal_samples[30281]=7021;
squeal_samples[30282]=4572;
squeal_samples[30283]=6461;
squeal_samples[30284]=9371;
squeal_samples[30285]=12150;
squeal_samples[30286]=14815;
squeal_samples[30287]=17357;
squeal_samples[30288]=19794;
squeal_samples[30289]=22115;
squeal_samples[30290]=24336;
squeal_samples[30291]=26463;
squeal_samples[30292]=28494;
squeal_samples[30293]=30429;
squeal_samples[30294]=32287;
squeal_samples[30295]=34055;
squeal_samples[30296]=35749;
squeal_samples[30297]=37358;
squeal_samples[30298]=38908;
squeal_samples[30299]=40374;
squeal_samples[30300]=41784;
squeal_samples[30301]=43127;
squeal_samples[30302]=44412;
squeal_samples[30303]=45637;
squeal_samples[30304]=46805;
squeal_samples[30305]=47927;
squeal_samples[30306]=48993;
squeal_samples[30307]=50012;
squeal_samples[30308]=50987;
squeal_samples[30309]=51919;
squeal_samples[30310]=52805;
squeal_samples[30311]=53654;
squeal_samples[30312]=54414;
squeal_samples[30313]=51042;
squeal_samples[30314]=45361;
squeal_samples[30315]=40052;
squeal_samples[30316]=35072;
squeal_samples[30317]=30424;
squeal_samples[30318]=26058;
squeal_samples[30319]=21985;
squeal_samples[30320]=18170;
squeal_samples[30321]=14599;
squeal_samples[30322]=11252;
squeal_samples[30323]=8128;
squeal_samples[30324]=5205;
squeal_samples[30325]=5322;
squeal_samples[30326]=8284;
squeal_samples[30327]=11113;
squeal_samples[30328]=13818;
squeal_samples[30329]=16411;
squeal_samples[30330]=18878;
squeal_samples[30331]=21243;
squeal_samples[30332]=23504;
squeal_samples[30333]=25666;
squeal_samples[30334]=27733;
squeal_samples[30335]=29702;
squeal_samples[30336]=31593;
squeal_samples[30337]=33392;
squeal_samples[30338]=35113;
squeal_samples[30339]=36752;
squeal_samples[30340]=38325;
squeal_samples[30341]=39822;
squeal_samples[30342]=41258;
squeal_samples[30343]=42618;
squeal_samples[30344]=43929;
squeal_samples[30345]=45170;
squeal_samples[30346]=46364;
squeal_samples[30347]=47500;
squeal_samples[30348]=48588;
squeal_samples[30349]=49624;
squeal_samples[30350]=50613;
squeal_samples[30351]=51560;
squeal_samples[30352]=52466;
squeal_samples[30353]=53333;
squeal_samples[30354]=54158;
squeal_samples[30355]=53039;
squeal_samples[30356]=47440;
squeal_samples[30357]=41986;
squeal_samples[30358]=36890;
squeal_samples[30359]=32115;
squeal_samples[30360]=27651;
squeal_samples[30361]=23472;
squeal_samples[30362]=19560;
squeal_samples[30363]=15895;
squeal_samples[30364]=12471;
squeal_samples[30365]=9261;
squeal_samples[30366]=6267;
squeal_samples[30367]=4582;
squeal_samples[30368]=7179;
squeal_samples[30369]=10053;
squeal_samples[30370]=12809;
squeal_samples[30371]=15436;
squeal_samples[30372]=17958;
squeal_samples[30373]=20355;
squeal_samples[30374]=22659;
squeal_samples[30375]=24855;
squeal_samples[30376]=26958;
squeal_samples[30377]=28963;
squeal_samples[30378]=30882;
squeal_samples[30379]=32713;
squeal_samples[30380]=34462;
squeal_samples[30381]=36134;
squeal_samples[30382]=37732;
squeal_samples[30383]=39260;
squeal_samples[30384]=40710;
squeal_samples[30385]=42103;
squeal_samples[30386]=43430;
squeal_samples[30387]=44701;
squeal_samples[30388]=45911;
squeal_samples[30389]=47066;
squeal_samples[30390]=48176;
squeal_samples[30391]=49226;
squeal_samples[30392]=50240;
squeal_samples[30393]=51198;
squeal_samples[30394]=52119;
squeal_samples[30395]=53001;
squeal_samples[30396]=53838;
squeal_samples[30397]=54168;
squeal_samples[30398]=49559;
squeal_samples[30399]=43984;
squeal_samples[30400]=38749;
squeal_samples[30401]=33860;
squeal_samples[30402]=29278;
squeal_samples[30403]=24993;
squeal_samples[30404]=20976;
squeal_samples[30405]=17233;
squeal_samples[30406]=13717;
squeal_samples[30407]=10431;
squeal_samples[30408]=7358;
squeal_samples[30409]=4657;
squeal_samples[30410]=6055;
squeal_samples[30411]=8975;
squeal_samples[30412]=11778;
squeal_samples[30413]=14453;
squeal_samples[30414]=17010;
squeal_samples[30415]=19463;
squeal_samples[30416]=21791;
squeal_samples[30417]=24034;
squeal_samples[30418]=26167;
squeal_samples[30419]=28213;
squeal_samples[30420]=30161;
squeal_samples[30421]=32026;
squeal_samples[30422]=33805;
squeal_samples[30423]=35507;
squeal_samples[30424]=37134;
squeal_samples[30425]=38679;
squeal_samples[30426]=40166;
squeal_samples[30427]=41580;
squeal_samples[30428]=42931;
squeal_samples[30429]=44223;
squeal_samples[30430]=45454;
squeal_samples[30431]=46633;
squeal_samples[30432]=47755;
squeal_samples[30433]=48827;
squeal_samples[30434]=49850;
squeal_samples[30435]=50838;
squeal_samples[30436]=51767;
squeal_samples[30437]=52666;
squeal_samples[30438]=53514;
squeal_samples[30439]=54339;
squeal_samples[30440]=51747;
squeal_samples[30441]=46016;
squeal_samples[30442]=40667;
squeal_samples[30443]=35639;
squeal_samples[30444]=30957;
squeal_samples[30445]=26551;
squeal_samples[30446]=22445;
squeal_samples[30447]=18600;
squeal_samples[30448]=14997;
squeal_samples[30449]=11628;
squeal_samples[30450]=8474;
squeal_samples[30451]=5525;
squeal_samples[30452]=4958;
squeal_samples[30453]=7885;
squeal_samples[30454]=10732;
squeal_samples[30455]=13454;
squeal_samples[30456]=16056;
squeal_samples[30457]=18547;
squeal_samples[30458]=20920;
squeal_samples[30459]=23195;
squeal_samples[30460]=25366;
squeal_samples[30461]=27444;
squeal_samples[30462]=29431;
squeal_samples[30463]=31325;
squeal_samples[30464]=33135;
squeal_samples[30465]=34870;
squeal_samples[30466]=36515;
squeal_samples[30467]=38099;
squeal_samples[30468]=39603;
squeal_samples[30469]=41044;
squeal_samples[30470]=42418;
squeal_samples[30471]=43737;
squeal_samples[30472]=44985;
squeal_samples[30473]=46185;
squeal_samples[30474]=47323;
squeal_samples[30475]=48420;
squeal_samples[30476]=49460;
squeal_samples[30477]=50459;
squeal_samples[30478]=51414;
squeal_samples[30479]=52316;
squeal_samples[30480]=53192;
squeal_samples[30481]=54024;
squeal_samples[30482]=53491;
squeal_samples[30483]=48111;
squeal_samples[30484]=42616;
squeal_samples[30485]=37476;
squeal_samples[30486]=32660;
squeal_samples[30487]=28164;
squeal_samples[30488]=23939;
squeal_samples[30489]=20002;
squeal_samples[30490]=16306;
squeal_samples[30491]=12854;
squeal_samples[30492]=9620;
squeal_samples[30493]=6597;
squeal_samples[30494]=4487;
squeal_samples[30495]=6778;
squeal_samples[30496]=9665;
squeal_samples[30497]=12432;
squeal_samples[30498]=15084;
squeal_samples[30499]=17612;
squeal_samples[30500]=20037;
squeal_samples[30501]=22340;
squeal_samples[30502]=24552;
squeal_samples[30503]=26667;
squeal_samples[30504]=28687;
squeal_samples[30505]=30614;
squeal_samples[30506]=32451;
squeal_samples[30507]=34218;
squeal_samples[30508]=35896;
squeal_samples[30509]=37507;
squeal_samples[30510]=39032;
squeal_samples[30511]=40501;
squeal_samples[30512]=41898;
squeal_samples[30513]=43235;
squeal_samples[30514]=44510;
squeal_samples[30515]=45729;
squeal_samples[30516]=46894;
squeal_samples[30517]=48002;
squeal_samples[30518]=49066;
squeal_samples[30519]=50077;
squeal_samples[30520]=51048;
squeal_samples[30521]=51974;
squeal_samples[30522]=52858;
squeal_samples[30523]=53700;
squeal_samples[30524]=54459;
squeal_samples[30525]=51074;
squeal_samples[30526]=45395;
squeal_samples[30527]=40073;
squeal_samples[30528]=35094;
squeal_samples[30529]=30439;
squeal_samples[30530]=26065;
squeal_samples[30531]=21991;
squeal_samples[30532]=18166;
squeal_samples[30533]=14598;
squeal_samples[30534]=11249;
squeal_samples[30535]=8121;
squeal_samples[30536]=5192;
squeal_samples[30537]=5310;
squeal_samples[30538]=8265;
squeal_samples[30539]=11094;
squeal_samples[30540]=13802;
squeal_samples[30541]=16383;
squeal_samples[30542]=18865;
squeal_samples[30543]=21214;
squeal_samples[30544]=23484;
squeal_samples[30545]=25640;
squeal_samples[30546]=27704;
squeal_samples[30547]=29674;
squeal_samples[30548]=31556;
squeal_samples[30549]=33359;
squeal_samples[30550]=35078;
squeal_samples[30551]=36718;
squeal_samples[30552]=38288;
squeal_samples[30553]=39791;
squeal_samples[30554]=41212;
squeal_samples[30555]=42585;
squeal_samples[30556]=43883;
squeal_samples[30557]=45133;
squeal_samples[30558]=46322;
squeal_samples[30559]=47460;
squeal_samples[30560]=48549;
squeal_samples[30561]=49581;
squeal_samples[30562]=50577;
squeal_samples[30563]=51513;
squeal_samples[30564]=52427;
squeal_samples[30565]=53282;
squeal_samples[30566]=54114;
squeal_samples[30567]=53574;
squeal_samples[30568]=48186;
squeal_samples[30569]=42686;
squeal_samples[30570]=37545;
squeal_samples[30571]=32719;
squeal_samples[30572]=28215;
squeal_samples[30573]=23989;
squeal_samples[30574]=20047;
squeal_samples[30575]=16350;
squeal_samples[30576]=12890;
squeal_samples[30577]=9651;
squeal_samples[30578]=6629;
squeal_samples[30579]=4512;
squeal_samples[30580]=6805;
squeal_samples[30581]=9684;
squeal_samples[30582]=12455;
squeal_samples[30583]=15096;
squeal_samples[30584]=17630;
squeal_samples[30585]=20049;
squeal_samples[30586]=22357;
squeal_samples[30587]=24566;
squeal_samples[30588]=26678;
squeal_samples[30589]=28691;
squeal_samples[30590]=30617;
squeal_samples[30591]=32463;
squeal_samples[30592]=34219;
squeal_samples[30593]=35899;
squeal_samples[30594]=37501;
squeal_samples[30595]=39041;
squeal_samples[30596]=40497;
squeal_samples[30597]=41898;
squeal_samples[30598]=43232;
squeal_samples[30599]=44509;
squeal_samples[30600]=45724;
squeal_samples[30601]=46891;
squeal_samples[30602]=47997;
squeal_samples[30603]=49057;
squeal_samples[30604]=50073;
squeal_samples[30605]=51038;
squeal_samples[30606]=51966;
squeal_samples[30607]=52848;
squeal_samples[30608]=53696;
squeal_samples[30609]=54451;
squeal_samples[30610]=51062;
squeal_samples[30611]=45383;
squeal_samples[30612]=40060;
squeal_samples[30613]=35085;
squeal_samples[30614]=30417;
squeal_samples[30615]=26057;
squeal_samples[30616]=21976;
squeal_samples[30617]=18155;
squeal_samples[30618]=14580;
squeal_samples[30619]=11232;
squeal_samples[30620]=8104;
squeal_samples[30621]=5172;
squeal_samples[30622]=5296;
squeal_samples[30623]=8245;
squeal_samples[30624]=11077;
squeal_samples[30625]=13785;
squeal_samples[30626]=16365;
squeal_samples[30627]=18841;
squeal_samples[30628]=21199;
squeal_samples[30629]=23458;
squeal_samples[30630]=25620;
squeal_samples[30631]=27684;
squeal_samples[30632]=29658;
squeal_samples[30633]=31538;
squeal_samples[30634]=33341;
squeal_samples[30635]=35056;
squeal_samples[30636]=36698;
squeal_samples[30637]=38268;
squeal_samples[30638]=39766;
squeal_samples[30639]=41196;
squeal_samples[30640]=42560;
squeal_samples[30641]=43867;
squeal_samples[30642]=45110;
squeal_samples[30643]=46303;
squeal_samples[30644]=47440;
squeal_samples[30645]=48521;
squeal_samples[30646]=49564;
squeal_samples[30647]=50549;
squeal_samples[30648]=51494;
squeal_samples[30649]=52400;
squeal_samples[30650]=53262;
squeal_samples[30651]=54088;
squeal_samples[30652]=53554;
squeal_samples[30653]=48166;
squeal_samples[30654]=42665;
squeal_samples[30655]=37519;
squeal_samples[30656]=32699;
squeal_samples[30657]=28190;
squeal_samples[30658]=23966;
squeal_samples[30659]=20026;
squeal_samples[30660]=16324;
squeal_samples[30661]=12869;
squeal_samples[30662]=9629;
squeal_samples[30663]=6602;
squeal_samples[30664]=4494;
squeal_samples[30665]=6777;
squeal_samples[30666]=9664;
squeal_samples[30667]=12430;
squeal_samples[30668]=15075;
squeal_samples[30669]=17605;
squeal_samples[30670]=20028;
squeal_samples[30671]=22332;
squeal_samples[30672]=24543;
squeal_samples[30673]=26657;
squeal_samples[30674]=28664;
squeal_samples[30675]=30598;
squeal_samples[30676]=32437;
squeal_samples[30677]=34198;
squeal_samples[30678]=35874;
squeal_samples[30679]=37480;
squeal_samples[30680]=39015;
squeal_samples[30681]=40476;
squeal_samples[30682]=41874;
squeal_samples[30683]=43211;
squeal_samples[30684]=44483;
squeal_samples[30685]=45703;
squeal_samples[30686]=46865;
squeal_samples[30687]=47977;
squeal_samples[30688]=49038;
squeal_samples[30689]=50050;
squeal_samples[30690]=51015;
squeal_samples[30691]=51942;
squeal_samples[30692]=52825;
squeal_samples[30693]=53674;
squeal_samples[30694]=54425;
squeal_samples[30695]=51042;
squeal_samples[30696]=45358;
squeal_samples[30697]=40038;
squeal_samples[30698]=35061;
squeal_samples[30699]=30394;
squeal_samples[30700]=26034;
squeal_samples[30701]=21953;
squeal_samples[30702]=18132;
squeal_samples[30703]=14556;
squeal_samples[30704]=11211;
squeal_samples[30705]=8078;
squeal_samples[30706]=5153;
squeal_samples[30707]=5268;
squeal_samples[30708]=8224;
squeal_samples[30709]=11054;
squeal_samples[30710]=13762;
squeal_samples[30711]=16342;
squeal_samples[30712]=18823;
squeal_samples[30713]=21174;
squeal_samples[30714]=23437;
squeal_samples[30715]=25596;
squeal_samples[30716]=27662;
squeal_samples[30717]=29633;
squeal_samples[30718]=31516;
squeal_samples[30719]=33317;
squeal_samples[30720]=35033;
squeal_samples[30721]=36676;
squeal_samples[30722]=38243;
squeal_samples[30723]=39744;
squeal_samples[30724]=41172;
squeal_samples[30725]=42537;
squeal_samples[30726]=43843;
squeal_samples[30727]=45087;
squeal_samples[30728]=46281;
squeal_samples[30729]=47414;
squeal_samples[30730]=48502;
squeal_samples[30731]=49536;
squeal_samples[30732]=50528;
squeal_samples[30733]=51472;
squeal_samples[30734]=52374;
squeal_samples[30735]=53242;
squeal_samples[30736]=54062;
squeal_samples[30737]=53532;
squeal_samples[30738]=48143;
squeal_samples[30739]=42641;
squeal_samples[30740]=37497;
squeal_samples[30741]=32675;
squeal_samples[30742]=28167;
squeal_samples[30743]=23944;
squeal_samples[30744]=19999;
squeal_samples[30745]=16305;
squeal_samples[30746]=12844;
squeal_samples[30747]=9606;
squeal_samples[30748]=6580;
squeal_samples[30749]=4467;
squeal_samples[30750]=6758;
squeal_samples[30751]=9637;
squeal_samples[30752]=12411;
squeal_samples[30753]=15047;
squeal_samples[30754]=17586;
squeal_samples[30755]=20000;
squeal_samples[30756]=22313;
squeal_samples[30757]=24518;
squeal_samples[30758]=26632;
squeal_samples[30759]=28644;
squeal_samples[30760]=30572;
squeal_samples[30761]=32414;
squeal_samples[30762]=34176;
squeal_samples[30763]=35848;
squeal_samples[30764]=37459;
squeal_samples[30765]=38991;
squeal_samples[30766]=40452;
squeal_samples[30767]=41851;
squeal_samples[30768]=43186;
squeal_samples[30769]=44463;
squeal_samples[30770]=45675;
squeal_samples[30771]=46847;
squeal_samples[30772]=47950;
squeal_samples[30773]=49015;
squeal_samples[30774]=50028;
squeal_samples[30775]=50990;
squeal_samples[30776]=51920;
squeal_samples[30777]=52802;
squeal_samples[30778]=53649;
squeal_samples[30779]=54403;
squeal_samples[30780]=51018;
squeal_samples[30781]=45334;
squeal_samples[30782]=40016;
squeal_samples[30783]=35036;
squeal_samples[30784]=30372;
squeal_samples[30785]=26010;
squeal_samples[30786]=21928;
squeal_samples[30787]=18111;
squeal_samples[30788]=14531;
squeal_samples[30789]=11187;
squeal_samples[30790]=8057;
squeal_samples[30791]=5125;
squeal_samples[30792]=5250;
squeal_samples[30793]=8197;
squeal_samples[30794]=11033;
squeal_samples[30795]=13735;
squeal_samples[30796]=16321;
squeal_samples[30797]=18799;
squeal_samples[30798]=21152;
squeal_samples[30799]=23412;
squeal_samples[30800]=25572;
squeal_samples[30801]=27639;
squeal_samples[30802]=29610;
squeal_samples[30803]=31493;
squeal_samples[30804]=33293;
squeal_samples[30805]=35009;
squeal_samples[30806]=36653;
squeal_samples[30807]=38219;
squeal_samples[30808]=39720;
squeal_samples[30809]=41151;
squeal_samples[30810]=42511;
squeal_samples[30811]=43822;
squeal_samples[30812]=45061;
squeal_samples[30813]=46259;
squeal_samples[30814]=47389;
squeal_samples[30815]=48481;
squeal_samples[30816]=49509;
squeal_samples[30817]=50508;
squeal_samples[30818]=51446;
squeal_samples[30819]=52351;
squeal_samples[30820]=53219;
squeal_samples[30821]=54037;
squeal_samples[30822]=53511;
squeal_samples[30823]=48116;
squeal_samples[30824]=42621;
squeal_samples[30825]=37470;
squeal_samples[30826]=32654;
squeal_samples[30827]=28142;
squeal_samples[30828]=23920;
squeal_samples[30829]=19978;
squeal_samples[30830]=16279;
squeal_samples[30831]=12821;
squeal_samples[30832]=9582;
squeal_samples[30833]=6556;
squeal_samples[30834]=4445;
squeal_samples[30835]=6734;
squeal_samples[30836]=9614;
squeal_samples[30837]=12386;
squeal_samples[30838]=15024;
squeal_samples[30839]=17561;
squeal_samples[30840]=19979;
squeal_samples[30841]=22287;
squeal_samples[30842]=24496;
squeal_samples[30843]=26608;
squeal_samples[30844]=28619;
squeal_samples[30845]=30550;
squeal_samples[30846]=32388;
squeal_samples[30847]=34155;
squeal_samples[30848]=35823;
squeal_samples[30849]=37436;
squeal_samples[30850]=38966;
squeal_samples[30851]=40429;
squeal_samples[30852]=41827;
squeal_samples[30853]=43165;
squeal_samples[30854]=44435;
squeal_samples[30855]=45656;
squeal_samples[30856]=46817;
squeal_samples[30857]=47931;
squeal_samples[30858]=48989;
squeal_samples[30859]=50005;
squeal_samples[30860]=50966;
squeal_samples[30861]=51895;
squeal_samples[30862]=52779;
squeal_samples[30863]=53623;
squeal_samples[30864]=54434;
squeal_samples[30865]=51824;
squeal_samples[30866]=46090;
squeal_samples[30867]=40717;
squeal_samples[30868]=35693;
squeal_samples[30869]=30987;
squeal_samples[30870]=26584;
squeal_samples[30871]=22460;
squeal_samples[30872]=18604;
squeal_samples[30873]=15001;
squeal_samples[30874]=11615;
squeal_samples[30875]=8466;
squeal_samples[30876]=5502;
squeal_samples[30877]=4937;
squeal_samples[30878]=7853;
squeal_samples[30879]=10698;
squeal_samples[30880]=13415;
squeal_samples[30881]=16013;
squeal_samples[30882]=18504;
squeal_samples[30883]=20874;
squeal_samples[30884]=23142;
squeal_samples[30885]=25316;
squeal_samples[30886]=27386;
squeal_samples[30887]=29371;
squeal_samples[30888]=31260;
squeal_samples[30889]=33078;
squeal_samples[30890]=34796;
squeal_samples[30891]=36454;
squeal_samples[30892]=38024;
squeal_samples[30893]=39536;
squeal_samples[30894]=40965;
squeal_samples[30895]=42346;
squeal_samples[30896]=43653;
squeal_samples[30897]=44904;
squeal_samples[30898]=46103;
squeal_samples[30899]=47241;
squeal_samples[30900]=48335;
squeal_samples[30901]=49375;
squeal_samples[30902]=50372;
squeal_samples[30903]=51320;
squeal_samples[30904]=52229;
squeal_samples[30905]=53099;
squeal_samples[30906]=53929;
squeal_samples[30907]=54243;
squeal_samples[30908]=49629;
squeal_samples[30909]=44032;
squeal_samples[30910]=38791;
squeal_samples[30911]=33886;
squeal_samples[30912]=29300;
squeal_samples[30913]=24995;
squeal_samples[30914]=20983;
squeal_samples[30915]=17218;
squeal_samples[30916]=13701;
squeal_samples[30917]=10405;
squeal_samples[30918]=7319;
squeal_samples[30919]=4620;
squeal_samples[30920]=6007;
squeal_samples[30921]=8933;
squeal_samples[30922]=11722;
squeal_samples[30923]=14396;
squeal_samples[30924]=16953;
squeal_samples[30925]=19397;
squeal_samples[30926]=21725;
squeal_samples[30927]=23962;
squeal_samples[30928]=26095;
squeal_samples[30929]=28135;
squeal_samples[30930]=30085;
squeal_samples[30931]=31944;
squeal_samples[30932]=33719;
squeal_samples[30933]=35419;
squeal_samples[30934]=37038;
squeal_samples[30935]=38594;
squeal_samples[30936]=40067;
squeal_samples[30937]=41482;
squeal_samples[30938]=42833;
squeal_samples[30939]=44117;
squeal_samples[30940]=45356;
squeal_samples[30941]=46523;
squeal_samples[30942]=47648;
squeal_samples[30943]=48725;
squeal_samples[30944]=49744;
squeal_samples[30945]=50722;
squeal_samples[30946]=51657;
squeal_samples[30947]=52548;
squeal_samples[30948]=53405;
squeal_samples[30949]=54222;
squeal_samples[30950]=53090;
squeal_samples[30951]=47475;
squeal_samples[30952]=42017;
squeal_samples[30953]=36904;
squeal_samples[30954]=32123;
squeal_samples[30955]=27638;
squeal_samples[30956]=23451;
squeal_samples[30957]=19533;
squeal_samples[30958]=15864;
squeal_samples[30959]=12426;
squeal_samples[30960]=9214;
squeal_samples[30961]=6205;
squeal_samples[30962]=4519;
squeal_samples[30963]=7108;
squeal_samples[30964]=9978;
squeal_samples[30965]=12727;
squeal_samples[30966]=15354;
squeal_samples[30967]=17873;
squeal_samples[30968]=20266;
squeal_samples[30969]=22569;
squeal_samples[30970]=24756;
squeal_samples[30971]=26861;
squeal_samples[30972]=28860;
squeal_samples[30973]=30779;
squeal_samples[30974]=32603;
squeal_samples[30975]=34356;
squeal_samples[30976]=36021;
squeal_samples[30977]=37623;
squeal_samples[30978]=39135;
squeal_samples[30979]=40596;
squeal_samples[30980]=41979;
squeal_samples[30981]=43313;
squeal_samples[30982]=44574;
squeal_samples[30983]=45787;
squeal_samples[30984]=46940;
squeal_samples[30985]=48046;
squeal_samples[30986]=49094;
squeal_samples[30987]=50110;
squeal_samples[30988]=51067;
squeal_samples[30989]=51988;
squeal_samples[30990]=52863;
squeal_samples[30991]=53703;
squeal_samples[30992]=54451;
squeal_samples[30993]=51061;
squeal_samples[30994]=45374;
squeal_samples[30995]=40045;
squeal_samples[30996]=35068;
squeal_samples[30997]=30388;
squeal_samples[30998]=26025;
squeal_samples[30999]=21931;
squeal_samples[31000]=18116;
squeal_samples[31001]=14533;
squeal_samples[31002]=11185;
squeal_samples[31003]=8052;
squeal_samples[31004]=5115;
squeal_samples[31005]=5235;
squeal_samples[31006]=8190;
squeal_samples[31007]=11014;
squeal_samples[31008]=13715;
squeal_samples[31009]=16299;
squeal_samples[31010]=18774;
squeal_samples[31011]=21133;
squeal_samples[31012]=23388;
squeal_samples[31013]=25546;
squeal_samples[31014]=27606;
squeal_samples[31015]=29576;
squeal_samples[31016]=31461;
squeal_samples[31017]=33259;
squeal_samples[31018]=34979;
squeal_samples[31019]=36617;
squeal_samples[31020]=38183;
squeal_samples[31021]=39681;
squeal_samples[31022]=41111;
squeal_samples[31023]=42475;
squeal_samples[31024]=43783;
squeal_samples[31025]=45023;
squeal_samples[31026]=46213;
squeal_samples[31027]=47350;
squeal_samples[31028]=48429;
squeal_samples[31029]=49476;
squeal_samples[31030]=50454;
squeal_samples[31031]=51409;
squeal_samples[31032]=52302;
squeal_samples[31033]=53172;
squeal_samples[31034]=53992;
squeal_samples[31035]=53939;
squeal_samples[31036]=48873;
squeal_samples[31037]=43324;
squeal_samples[31038]=38122;
squeal_samples[31039]=33267;
squeal_samples[31040]=28706;
squeal_samples[31041]=24448;
squeal_samples[31042]=20458;
squeal_samples[31043]=16732;
squeal_samples[31044]=13235;
squeal_samples[31045]=9976;
squeal_samples[31046]=6912;
squeal_samples[31047]=4463;
squeal_samples[31048]=6344;
squeal_samples[31049]=9248;
squeal_samples[31050]=12028;
squeal_samples[31051]=14687;
squeal_samples[31052]=17224;
squeal_samples[31053]=19661;
squeal_samples[31054]=21977;
squeal_samples[31055]=24196;
squeal_samples[31056]=26321;
squeal_samples[31057]=28348;
squeal_samples[31058]=30280;
squeal_samples[31059]=32133;
squeal_samples[31060]=33898;
squeal_samples[31061]=35590;
squeal_samples[31062]=37204;
squeal_samples[31063]=38739;
squeal_samples[31064]=40211;
squeal_samples[31065]=41615;
squeal_samples[31066]=42962;
squeal_samples[31067]=44243;
squeal_samples[31068]=45462;
squeal_samples[31069]=46635;
squeal_samples[31070]=47748;
squeal_samples[31071]=48817;
squeal_samples[31072]=49834;
squeal_samples[31073]=50805;
squeal_samples[31074]=51736;
squeal_samples[31075]=52619;
squeal_samples[31076]=53473;
squeal_samples[31077]=54283;
squeal_samples[31078]=52468;
squeal_samples[31079]=46739;
squeal_samples[31080]=41321;
squeal_samples[31081]=36251;
squeal_samples[31082]=31509;
squeal_samples[31083]=27066;
squeal_samples[31084]=22910;
squeal_samples[31085]=19023;
squeal_samples[31086]=15383;
squeal_samples[31087]=11976;
squeal_samples[31088]=8788;
squeal_samples[31089]=5810;
squeal_samples[31090]=4633;
squeal_samples[31091]=7438;
squeal_samples[31092]=10293;
squeal_samples[31093]=13028;
squeal_samples[31094]=15640;
squeal_samples[31095]=18143;
squeal_samples[31096]=20527;
squeal_samples[31097]=22811;
squeal_samples[31098]=24994;
squeal_samples[31099]=27077;
squeal_samples[31100]=29071;
squeal_samples[31101]=30973;
squeal_samples[31102]=32793;
squeal_samples[31103]=34532;
squeal_samples[31104]=36191;
squeal_samples[31105]=37770;
squeal_samples[31106]=39295;
squeal_samples[31107]=40733;
squeal_samples[31108]=42115;
squeal_samples[31109]=43437;
squeal_samples[31110]=44697;
squeal_samples[31111]=45895;
squeal_samples[31112]=47048;
squeal_samples[31113]=48141;
squeal_samples[31114]=49192;
squeal_samples[31115]=50190;
squeal_samples[31116]=51147;
squeal_samples[31117]=52059;
squeal_samples[31118]=52933;
squeal_samples[31119]=53765;
squeal_samples[31120]=54355;
squeal_samples[31121]=50294;
squeal_samples[31122]=44652;
squeal_samples[31123]=39371;
squeal_samples[31124]=34424;
squeal_samples[31125]=29796;
squeal_samples[31126]=25466;
squeal_samples[31127]=21406;
squeal_samples[31128]=17619;
squeal_samples[31129]=14066;
squeal_samples[31130]=10741;
squeal_samples[31131]=7636;
squeal_samples[31132]=4775;
squeal_samples[31133]=5573;
squeal_samples[31134]=8514;
squeal_samples[31135]=11316;
squeal_samples[31136]=14013;
squeal_samples[31137]=16577;
squeal_samples[31138]=19037;
squeal_samples[31139]=21383;
squeal_samples[31140]=23630;
squeal_samples[31141]=25773;
squeal_samples[31142]=27827;
squeal_samples[31143]=29783;
squeal_samples[31144]=31657;
squeal_samples[31145]=33442;
squeal_samples[31146]=35150;
squeal_samples[31147]=36780;
squeal_samples[31148]=38339;
squeal_samples[31149]=39831;
squeal_samples[31150]=41246;
squeal_samples[31151]=42610;
squeal_samples[31152]=43899;
squeal_samples[31153]=45143;
squeal_samples[31154]=46321;
squeal_samples[31155]=47453;
squeal_samples[31156]=48528;
squeal_samples[31157]=49557;
squeal_samples[31158]=50543;
squeal_samples[31159]=51481;
squeal_samples[31160]=52380;
squeal_samples[31161]=53239;
squeal_samples[31162]=54059;
squeal_samples[31163]=53517;
squeal_samples[31164]=48121;
squeal_samples[31165]=42620;
squeal_samples[31166]=37460;
squeal_samples[31167]=32645;
squeal_samples[31168]=28120;
squeal_samples[31169]=23900;
squeal_samples[31170]=19945;
squeal_samples[31171]=16248;
squeal_samples[31172]=12782;
squeal_samples[31173]=9541;
squeal_samples[31174]=6511;
squeal_samples[31175]=4801;
squeal_samples[31176]=7372;
squeal_samples[31177]=10232;
squeal_samples[31178]=12965;
squeal_samples[31179]=15581;
squeal_samples[31180]=18088;
squeal_samples[31181]=20466;
squeal_samples[31182]=22758;
squeal_samples[31183]=24939;
squeal_samples[31184]=27027;
squeal_samples[31185]=29024;
squeal_samples[31186]=30925;
squeal_samples[31187]=32750;
squeal_samples[31188]=34478;
squeal_samples[31189]=36145;
squeal_samples[31190]=37731;
squeal_samples[31191]=39246;
squeal_samples[31192]=40694;
squeal_samples[31193]=42074;
squeal_samples[31194]=43390;
squeal_samples[31195]=44657;
squeal_samples[31196]=45854;
squeal_samples[31197]=47006;
squeal_samples[31198]=48101;
squeal_samples[31199]=49152;
squeal_samples[31200]=50153;
squeal_samples[31201]=51111;
squeal_samples[31202]=52026;
squeal_samples[31203]=52892;
squeal_samples[31204]=53737;
squeal_samples[31205]=54475;
squeal_samples[31206]=51088;
squeal_samples[31207]=45387;
squeal_samples[31208]=40058;
squeal_samples[31209]=35068;
squeal_samples[31210]=30396;
squeal_samples[31211]=26022;
squeal_samples[31212]=21930;
squeal_samples[31213]=18105;
squeal_samples[31214]=14518;
squeal_samples[31215]=11170;
squeal_samples[31216]=8033;
squeal_samples[31217]=5099;
squeal_samples[31218]=5212;
squeal_samples[31219]=8161;
squeal_samples[31220]=10985;
squeal_samples[31221]=13687;
squeal_samples[31222]=16271;
squeal_samples[31223]=18741;
squeal_samples[31224]=21099;
squeal_samples[31225]=23353;
squeal_samples[31226]=25513;
squeal_samples[31227]=27573;
squeal_samples[31228]=29542;
squeal_samples[31229]=31427;
squeal_samples[31230]=33221;
squeal_samples[31231]=34936;
squeal_samples[31232]=36576;
squeal_samples[31233]=38144;
squeal_samples[31234]=39639;
squeal_samples[31235]=41069;
squeal_samples[31236]=42429;
squeal_samples[31237]=43731;
squeal_samples[31238]=44982;
squeal_samples[31239]=46167;
squeal_samples[31240]=47303;
squeal_samples[31241]=48384;
squeal_samples[31242]=49419;
squeal_samples[31243]=50410;
squeal_samples[31244]=51352;
squeal_samples[31245]=52260;
squeal_samples[31246]=53114;
squeal_samples[31247]=53946;
squeal_samples[31248]=54256;
squeal_samples[31249]=49625;
squeal_samples[31250]=44033;
squeal_samples[31251]=38776;
squeal_samples[31252]=33874;
squeal_samples[31253]=29276;
squeal_samples[31254]=24976;
squeal_samples[31255]=20949;
squeal_samples[31256]=17183;
squeal_samples[31257]=13662;
squeal_samples[31258]=10361;
squeal_samples[31259]=7279;
squeal_samples[31260]=4568;
squeal_samples[31261]=5957;
squeal_samples[31262]=8876;
squeal_samples[31263]=11670;
squeal_samples[31264]=14340;
squeal_samples[31265]=16897;
squeal_samples[31266]=19334;
squeal_samples[31267]=21669;
squeal_samples[31268]=23895;
squeal_samples[31269]=26032;
squeal_samples[31270]=28064;
squeal_samples[31271]=30015;
squeal_samples[31272]=31874;
squeal_samples[31273]=33648;
squeal_samples[31274]=35350;
squeal_samples[31275]=36968;
squeal_samples[31276]=38518;
squeal_samples[31277]=39991;
squeal_samples[31278]=41406;
squeal_samples[31279]=42757;
squeal_samples[31280]=44037;
squeal_samples[31281]=45275;
squeal_samples[31282]=46441;
squeal_samples[31283]=47569;
squeal_samples[31284]=48635;
squeal_samples[31285]=49665;
squeal_samples[31286]=50639;
squeal_samples[31287]=51578;
squeal_samples[31288]=52466;
squeal_samples[31289]=53317;
squeal_samples[31290]=54136;
squeal_samples[31291]=53582;
squeal_samples[31292]=48191;
squeal_samples[31293]=42672;
squeal_samples[31294]=37513;
squeal_samples[31295]=32689;
squeal_samples[31296]=28158;
squeal_samples[31297]=23936;
squeal_samples[31298]=19979;
squeal_samples[31299]=16270;
squeal_samples[31300]=12807;
squeal_samples[31301]=9558;
squeal_samples[31302]=6524;
squeal_samples[31303]=4408;
squeal_samples[31304]=6686;
squeal_samples[31305]=9579;
squeal_samples[31306]=12335;
squeal_samples[31307]=14975;
squeal_samples[31308]=17509;
squeal_samples[31309]=19913;
squeal_samples[31310]=22229;
squeal_samples[31311]=24422;
squeal_samples[31312]=26545;
squeal_samples[31313]=28547;
squeal_samples[31314]=30477;
squeal_samples[31315]=32313;
squeal_samples[31316]=34067;
squeal_samples[31317]=35754;
squeal_samples[31318]=37342;
squeal_samples[31319]=38883;
squeal_samples[31320]=40340;
squeal_samples[31321]=41740;
squeal_samples[31322]=43070;
squeal_samples[31323]=44345;
squeal_samples[31324]=45555;
squeal_samples[31325]=46721;
squeal_samples[31326]=47826;
squeal_samples[31327]=48885;
squeal_samples[31328]=49902;
squeal_samples[31329]=50866;
squeal_samples[31330]=51788;
squeal_samples[31331]=52671;
squeal_samples[31332]=53514;
squeal_samples[31333]=54318;
squeal_samples[31334]=52503;
squeal_samples[31335]=46763;
squeal_samples[31336]=41340;
squeal_samples[31337]=36265;
squeal_samples[31338]=31510;
squeal_samples[31339]=27071;
squeal_samples[31340]=22904;
squeal_samples[31341]=19018;
squeal_samples[31342]=15372;
squeal_samples[31343]=11965;
squeal_samples[31344]=8766;
squeal_samples[31345]=5788;
squeal_samples[31346]=4607;
squeal_samples[31347]=7414;
squeal_samples[31348]=10264;
squeal_samples[31349]=12996;
squeal_samples[31350]=15613;
squeal_samples[31351]=18104;
squeal_samples[31352]=20493;
squeal_samples[31353]=22771;
squeal_samples[31354]=24952;
squeal_samples[31355]=27039;
squeal_samples[31356]=29026;
squeal_samples[31357]=30930;
squeal_samples[31358]=32744;
squeal_samples[31359]=34484;
squeal_samples[31360]=36140;
squeal_samples[31361]=37729;
squeal_samples[31362]=39239;
squeal_samples[31363]=40684;
squeal_samples[31364]=42063;
squeal_samples[31365]=43377;
squeal_samples[31366]=44644;
squeal_samples[31367]=45840;
squeal_samples[31368]=46993;
squeal_samples[31369]=48082;
squeal_samples[31370]=49137;
squeal_samples[31371]=50130;
squeal_samples[31372]=51093;
squeal_samples[31373]=51998;
squeal_samples[31374]=52877;
squeal_samples[31375]=53704;
squeal_samples[31376]=54452;
squeal_samples[31377]=51053;
squeal_samples[31378]=45361;
squeal_samples[31379]=40025;
squeal_samples[31380]=35035;
squeal_samples[31381]=30364;
squeal_samples[31382]=25988;
squeal_samples[31383]=21893;
squeal_samples[31384]=18073;
squeal_samples[31385]=14484;
squeal_samples[31386]=11134;
squeal_samples[31387]=7992;
squeal_samples[31388]=5063;
squeal_samples[31389]=5167;
squeal_samples[31390]=8124;
squeal_samples[31391]=10947;
squeal_samples[31392]=13649;
squeal_samples[31393]=16231;
squeal_samples[31394]=18700;
squeal_samples[31395]=21053;
squeal_samples[31396]=23313;
squeal_samples[31397]=25472;
squeal_samples[31398]=27530;
squeal_samples[31399]=29498;
squeal_samples[31400]=31385;
squeal_samples[31401]=33175;
squeal_samples[31402]=34896;
squeal_samples[31403]=36530;
squeal_samples[31404]=38100;
squeal_samples[31405]=39592;
squeal_samples[31406]=41023;
squeal_samples[31407]=42387;
squeal_samples[31408]=43688;
squeal_samples[31409]=44930;
squeal_samples[31410]=46122;
squeal_samples[31411]=47250;
squeal_samples[31412]=48344;
squeal_samples[31413]=49372;
squeal_samples[31414]=50369;
squeal_samples[31415]=51303;
squeal_samples[31416]=52208;
squeal_samples[31417]=53074;
squeal_samples[31418]=53895;
squeal_samples[31419]=54206;
squeal_samples[31420]=49586;
squeal_samples[31421]=43977;
squeal_samples[31422]=38740;
squeal_samples[31423]=33823;
squeal_samples[31424]=29232;
squeal_samples[31425]=24925;
squeal_samples[31426]=20900;
squeal_samples[31427]=17141;
squeal_samples[31428]=13611;
squeal_samples[31429]=10313;
squeal_samples[31430]=7230;
squeal_samples[31431]=4518;
squeal_samples[31432]=5910;
squeal_samples[31433]=8827;
squeal_samples[31434]=11620;
squeal_samples[31435]=14292;
squeal_samples[31436]=16846;
squeal_samples[31437]=19288;
squeal_samples[31438]=21618;
squeal_samples[31439]=23849;
squeal_samples[31440]=25979;
squeal_samples[31441]=28018;
squeal_samples[31442]=29964;
squeal_samples[31443]=31826;
squeal_samples[31444]=33601;
squeal_samples[31445]=35298;
squeal_samples[31446]=36919;
squeal_samples[31447]=38470;
squeal_samples[31448]=39941;
squeal_samples[31449]=41360;
squeal_samples[31450]=42705;
squeal_samples[31451]=43994;
squeal_samples[31452]=45225;
squeal_samples[31453]=46398;
squeal_samples[31454]=47520;
squeal_samples[31455]=48592;
squeal_samples[31456]=49615;
squeal_samples[31457]=50592;
squeal_samples[31458]=51525;
squeal_samples[31459]=52421;
squeal_samples[31460]=53265;
squeal_samples[31461]=54089;
squeal_samples[31462]=53533;
squeal_samples[31463]=48141;
squeal_samples[31464]=42623;
squeal_samples[31465]=37466;
squeal_samples[31466]=32635;
squeal_samples[31467]=28115;
squeal_samples[31468]=23882;
squeal_samples[31469]=19932;
squeal_samples[31470]=16220;
squeal_samples[31471]=12757;
squeal_samples[31472]=9514;
squeal_samples[31473]=6475;
squeal_samples[31474]=4765;
squeal_samples[31475]=7333;
squeal_samples[31476]=10192;
squeal_samples[31477]=12920;
squeal_samples[31478]=15542;
squeal_samples[31479]=18037;
squeal_samples[31480]=20422;
squeal_samples[31481]=22706;
squeal_samples[31482]=24890;
squeal_samples[31483]=26971;
squeal_samples[31484]=28966;
squeal_samples[31485]=30869;
squeal_samples[31486]=32687;
squeal_samples[31487]=34424;
squeal_samples[31488]=36083;
squeal_samples[31489]=37667;
squeal_samples[31490]=39184;
squeal_samples[31491]=40629;
squeal_samples[31492]=42009;
squeal_samples[31493]=43328;
squeal_samples[31494]=44585;
squeal_samples[31495]=45792;
squeal_samples[31496]=46936;
squeal_samples[31497]=48037;
squeal_samples[31498]=49081;
squeal_samples[31499]=50086;
squeal_samples[31500]=51040;
squeal_samples[31501]=51957;
squeal_samples[31502]=52822;
squeal_samples[31503]=53660;
squeal_samples[31504]=54456;
squeal_samples[31505]=51844;
squeal_samples[31506]=46095;
squeal_samples[31507]=40710;
squeal_samples[31508]=35672;
squeal_samples[31509]=30957;
squeal_samples[31510]=26543;
squeal_samples[31511]=22411;
squeal_samples[31512]=18550;
squeal_samples[31513]=14934;
squeal_samples[31514]=11544;
squeal_samples[31515]=8378;
squeal_samples[31516]=5413;
squeal_samples[31517]=4841;
squeal_samples[31518]=7758;
squeal_samples[31519]=10597;
squeal_samples[31520]=13312;
squeal_samples[31521]=15908;
squeal_samples[31522]=18391;
squeal_samples[31523]=20755;
squeal_samples[31524]=23028;
squeal_samples[31525]=25195;
squeal_samples[31526]=27267;
squeal_samples[31527]=29243;
squeal_samples[31528]=31136;
squeal_samples[31529]=32941;
squeal_samples[31530]=34665;
squeal_samples[31531]=36318;
squeal_samples[31532]=37886;
squeal_samples[31533]=39396;
squeal_samples[31534]=40827;
squeal_samples[31535]=42200;
squeal_samples[31536]=43509;
squeal_samples[31537]=44758;
squeal_samples[31538]=45954;
squeal_samples[31539]=47091;
squeal_samples[31540]=48184;
squeal_samples[31541]=49225;
squeal_samples[31542]=50221;
squeal_samples[31543]=51163;
squeal_samples[31544]=52075;
squeal_samples[31545]=52936;
squeal_samples[31546]=53767;
squeal_samples[31547]=54511;
squeal_samples[31548]=51107;
squeal_samples[31549]=45405;
squeal_samples[31550]=40061;
squeal_samples[31551]=35069;
squeal_samples[31552]=30391;
squeal_samples[31553]=26009;
squeal_samples[31554]=21916;
squeal_samples[31555]=18082;
squeal_samples[31556]=14497;
squeal_samples[31557]=11136;
squeal_samples[31558]=7995;
squeal_samples[31559]=5055;
squeal_samples[31560]=5171;
squeal_samples[31561]=8115;
squeal_samples[31562]=10937;
squeal_samples[31563]=13638;
squeal_samples[31564]=16220;
squeal_samples[31565]=18691;
squeal_samples[31566]=21040;
squeal_samples[31567]=23297;
squeal_samples[31568]=25451;
squeal_samples[31569]=27512;
squeal_samples[31570]=29479;
squeal_samples[31571]=31359;
squeal_samples[31572]=33158;
squeal_samples[31573]=34870;
squeal_samples[31574]=36511;
squeal_samples[31575]=38072;
squeal_samples[31576]=39569;
squeal_samples[31577]=40998;
squeal_samples[31578]=42358;
squeal_samples[31579]=43662;
squeal_samples[31580]=44904;
squeal_samples[31581]=46091;
squeal_samples[31582]=47228;
squeal_samples[31583]=48305;
squeal_samples[31584]=49346;
squeal_samples[31585]=50325;
squeal_samples[31586]=51274;
squeal_samples[31587]=52174;
squeal_samples[31588]=53035;
squeal_samples[31589]=53858;
squeal_samples[31590]=54432;
squeal_samples[31591]=50364;
squeal_samples[31592]=44705;
squeal_samples[31593]=39412;
squeal_samples[31594]=34456;
squeal_samples[31595]=29815;
squeal_samples[31596]=25477;
squeal_samples[31597]=21407;
squeal_samples[31598]=17615;
squeal_samples[31599]=14051;
squeal_samples[31600]=10721;
squeal_samples[31601]=7610;
squeal_samples[31602]=4736;
squeal_samples[31603]=5533;
squeal_samples[31604]=8465;
squeal_samples[31605]=11271;
squeal_samples[31606]=13957;
squeal_samples[31607]=16524;
squeal_samples[31608]=18979;
squeal_samples[31609]=21320;
squeal_samples[31610]=23560;
squeal_samples[31611]=25704;
squeal_samples[31612]=27752;
squeal_samples[31613]=29708;
squeal_samples[31614]=31577;
squeal_samples[31615]=33362;
squeal_samples[31616]=35064;
squeal_samples[31617]=36701;
squeal_samples[31618]=38248;
squeal_samples[31619]=39738;
squeal_samples[31620]=41158;
squeal_samples[31621]=42514;
squeal_samples[31622]=43809;
squeal_samples[31623]=45041;
squeal_samples[31624]=46222;
squeal_samples[31625]=47351;
squeal_samples[31626]=48423;
squeal_samples[31627]=49460;
squeal_samples[31628]=50437;
squeal_samples[31629]=51375;
squeal_samples[31630]=52273;
squeal_samples[31631]=53129;
squeal_samples[31632]=53952;
squeal_samples[31633]=54251;
squeal_samples[31634]=49623;
squeal_samples[31635]=44016;
squeal_samples[31636]=38761;
squeal_samples[31637]=33851;
squeal_samples[31638]=29240;
squeal_samples[31639]=24940;
squeal_samples[31640]=20906;
squeal_samples[31641]=17141;
squeal_samples[31642]=13610;
squeal_samples[31643]=10307;
squeal_samples[31644]=7223;
squeal_samples[31645]=4506;
squeal_samples[31646]=5898;
squeal_samples[31647]=8807;
squeal_samples[31648]=11606;
squeal_samples[31649]=14268;
squeal_samples[31650]=16823;
squeal_samples[31651]=19266;
squeal_samples[31652]=21593;
squeal_samples[31653]=23821;
squeal_samples[31654]=25952;
squeal_samples[31655]=27989;
squeal_samples[31656]=29936;
squeal_samples[31657]=31793;
squeal_samples[31658]=33565;
squeal_samples[31659]=35266;
squeal_samples[31660]=36880;
squeal_samples[31661]=38430;
squeal_samples[31662]=39907;
squeal_samples[31663]=41323;
squeal_samples[31664]=42662;
squeal_samples[31665]=43955;
squeal_samples[31666]=45181;
squeal_samples[31667]=46357;
squeal_samples[31668]=47472;
squeal_samples[31669]=48551;
squeal_samples[31670]=49567;
squeal_samples[31671]=50551;
squeal_samples[31672]=51473;
squeal_samples[31673]=52369;
squeal_samples[31674]=53224;
squeal_samples[31675]=54033;
squeal_samples[31676]=53968;
squeal_samples[31677]=48889;
squeal_samples[31678]=43327;
squeal_samples[31679]=38119;
squeal_samples[31680]=33245;
squeal_samples[31681]=28676;
squeal_samples[31682]=24410;
squeal_samples[31683]=20412;
squeal_samples[31684]=16678;
squeal_samples[31685]=13174;
squeal_samples[31686]=9899;
squeal_samples[31687]=6834;
squeal_samples[31688]=4377;
squeal_samples[31689]=6251;
squeal_samples[31690]=9160;
squeal_samples[31691]=11925;
squeal_samples[31692]=14586;
squeal_samples[31693]=17123;
squeal_samples[31694]=19553;
squeal_samples[31695]=21863;
squeal_samples[31696]=24082;
squeal_samples[31697]=26199;
squeal_samples[31698]=28227;
squeal_samples[31699]=30157;
squeal_samples[31700]=32008;
squeal_samples[31701]=33771;
squeal_samples[31702]=35460;
squeal_samples[31703]=37069;
squeal_samples[31704]=38606;
squeal_samples[31705]=40077;
squeal_samples[31706]=41475;
squeal_samples[31707]=42817;
squeal_samples[31708]=44096;
squeal_samples[31709]=45318;
squeal_samples[31710]=46485;
squeal_samples[31711]=47603;
squeal_samples[31712]=48666;
squeal_samples[31713]=49683;
squeal_samples[31714]=50655;
squeal_samples[31715]=51577;
squeal_samples[31716]=52467;
squeal_samples[31717]=53312;
squeal_samples[31718]=54124;
squeal_samples[31719]=53570;
squeal_samples[31720]=48164;
squeal_samples[31721]=42644;
squeal_samples[31722]=37477;
squeal_samples[31723]=32649;
squeal_samples[31724]=28112;
squeal_samples[31725]=23886;
squeal_samples[31726]=19918;
squeal_samples[31727]=16219;
squeal_samples[31728]=12740;
squeal_samples[31729]=9499;
squeal_samples[31730]=6450;
squeal_samples[31731]=4333;
squeal_samples[31732]=6611;
squeal_samples[31733]=9498;
squeal_samples[31734]=12257;
squeal_samples[31735]=14899;
squeal_samples[31736]=17420;
squeal_samples[31737]=19836;
squeal_samples[31738]=22131;
squeal_samples[31739]=24343;
squeal_samples[31740]=26440;
squeal_samples[31741]=28462;
squeal_samples[31742]=30380;
squeal_samples[31743]=32221;
squeal_samples[31744]=33975;
squeal_samples[31745]=35654;
squeal_samples[31746]=37253;
squeal_samples[31747]=38784;
squeal_samples[31748]=40242;
squeal_samples[31749]=41638;
squeal_samples[31750]=42968;
squeal_samples[31751]=44241;
squeal_samples[31752]=45458;
squeal_samples[31753]=46614;
squeal_samples[31754]=47725;
squeal_samples[31755]=48782;
squeal_samples[31756]=49792;
squeal_samples[31757]=50760;
squeal_samples[31758]=51678;
squeal_samples[31759]=52564;
squeal_samples[31760]=53402;
squeal_samples[31761]=54211;
squeal_samples[31762]=53068;
squeal_samples[31763]=47442;
squeal_samples[31764]=41968;
squeal_samples[31765]=36846;
squeal_samples[31766]=32053;
squeal_samples[31767]=27562;
squeal_samples[31768]=23357;
squeal_samples[31769]=19435;
squeal_samples[31770]=15748;
squeal_samples[31771]=12316;
squeal_samples[31772]=9089;
squeal_samples[31773]=6079;
squeal_samples[31774]=4870;
squeal_samples[31775]=7662;
squeal_samples[31776]=10492;
squeal_samples[31777]=13216;
squeal_samples[31778]=15810;
squeal_samples[31779]=18299;
squeal_samples[31780]=20658;
squeal_samples[31781]=22935;
squeal_samples[31782]=25099;
squeal_samples[31783]=27178;
squeal_samples[31784]=29156;
squeal_samples[31785]=31044;
squeal_samples[31786]=32854;
squeal_samples[31787]=34574;
squeal_samples[31788]=36230;
squeal_samples[31789]=37798;
squeal_samples[31790]=39310;
squeal_samples[31791]=40741;
squeal_samples[31792]=42112;
squeal_samples[31793]=43424;
squeal_samples[31794]=44673;
squeal_samples[31795]=45870;
squeal_samples[31796]=47009;
squeal_samples[31797]=48098;
squeal_samples[31798]=49145;
squeal_samples[31799]=50133;
squeal_samples[31800]=51090;
squeal_samples[31801]=51992;
squeal_samples[31802]=52861;
squeal_samples[31803]=53690;
squeal_samples[31804]=54423;
squeal_samples[31805]=51034;
squeal_samples[31806]=45322;
squeal_samples[31807]=39986;
squeal_samples[31808]=34990;
squeal_samples[31809]=30313;
squeal_samples[31810]=25936;
squeal_samples[31811]=21838;
squeal_samples[31812]=18007;
squeal_samples[31813]=14421;
squeal_samples[31814]=11063;
squeal_samples[31815]=7916;
squeal_samples[31816]=5026;
squeal_samples[31817]=5801;
squeal_samples[31818]=8724;
squeal_samples[31819]=11516;
squeal_samples[31820]=14183;
squeal_samples[31821]=16742;
squeal_samples[31822]=19184;
squeal_samples[31823]=21513;
squeal_samples[31824]=23744;
squeal_samples[31825]=25878;
squeal_samples[31826]=27912;
squeal_samples[31827]=29863;
squeal_samples[31828]=31714;
squeal_samples[31829]=33498;
squeal_samples[31830]=35188;
squeal_samples[31831]=36813;
squeal_samples[31832]=38358;
squeal_samples[31833]=39838;
squeal_samples[31834]=41251;
squeal_samples[31835]=42600;
squeal_samples[31836]=43889;
squeal_samples[31837]=45111;
squeal_samples[31838]=46293;
squeal_samples[31839]=47413;
squeal_samples[31840]=48485;
squeal_samples[31841]=49505;
squeal_samples[31842]=50482;
squeal_samples[31843]=51418;
squeal_samples[31844]=52309;
squeal_samples[31845]=53161;
squeal_samples[31846]=53980;
squeal_samples[31847]=54268;
squeal_samples[31848]=49651;
squeal_samples[31849]=44019;
squeal_samples[31850]=38777;
squeal_samples[31851]=33851;
squeal_samples[31852]=29249;
squeal_samples[31853]=24936;
squeal_samples[31854]=20903;
squeal_samples[31855]=17127;
squeal_samples[31856]=13601;
squeal_samples[31857]=10288;
squeal_samples[31858]=7203;
squeal_samples[31859]=4482;
squeal_samples[31860]=5871;
squeal_samples[31861]=8786;
squeal_samples[31862]=11576;
squeal_samples[31863]=14242;
squeal_samples[31864]=16795;
squeal_samples[31865]=19231;
squeal_samples[31866]=21563;
squeal_samples[31867]=23786;
squeal_samples[31868]=25919;
squeal_samples[31869]=27957;
squeal_samples[31870]=29896;
squeal_samples[31871]=31755;
squeal_samples[31872]=33528;
squeal_samples[31873]=35219;
squeal_samples[31874]=36846;
squeal_samples[31875]=38387;
squeal_samples[31876]=39868;
squeal_samples[31877]=41274;
squeal_samples[31878]=42622;
squeal_samples[31879]=43909;
squeal_samples[31880]=45133;
squeal_samples[31881]=46307;
squeal_samples[31882]=47429;
squeal_samples[31883]=48500;
squeal_samples[31884]=49519;
squeal_samples[31885]=50500;
squeal_samples[31886]=51424;
squeal_samples[31887]=52322;
squeal_samples[31888]=53170;
squeal_samples[31889]=53988;
squeal_samples[31890]=54282;
squeal_samples[31891]=49648;
squeal_samples[31892]=44036;
squeal_samples[31893]=38777;
squeal_samples[31894]=33858;
squeal_samples[31895]=29245;
squeal_samples[31896]=24938;
squeal_samples[31897]=20898;
squeal_samples[31898]=17136;
squeal_samples[31899]=13595;
squeal_samples[31900]=10291;
squeal_samples[31901]=7197;
squeal_samples[31902]=4486;
squeal_samples[31903]=5865;
squeal_samples[31904]=8784;
squeal_samples[31905]=11566;
squeal_samples[31906]=14237;
squeal_samples[31907]=16788;
squeal_samples[31908]=19225;
squeal_samples[31909]=21557;
squeal_samples[31910]=23777;
squeal_samples[31911]=25916;
squeal_samples[31912]=27947;
squeal_samples[31913]=29893;
squeal_samples[31914]=31746;
squeal_samples[31915]=33521;
squeal_samples[31916]=35215;
squeal_samples[31917]=36836;
squeal_samples[31918]=38379;
squeal_samples[31919]=39858;
squeal_samples[31920]=41264;
squeal_samples[31921]=42615;
squeal_samples[31922]=43902;
squeal_samples[31923]=45125;
squeal_samples[31924]=46303;
squeal_samples[31925]=47415;
squeal_samples[31926]=48489;
squeal_samples[31927]=49513;
squeal_samples[31928]=50486;
squeal_samples[31929]=51420;
squeal_samples[31930]=52313;
squeal_samples[31931]=53159;
squeal_samples[31932]=53977;
squeal_samples[31933]=54269;
squeal_samples[31934]=49643;
squeal_samples[31935]=44023;
squeal_samples[31936]=38764;
squeal_samples[31937]=33847;
squeal_samples[31938]=29240;
squeal_samples[31939]=24928;
squeal_samples[31940]=20891;
squeal_samples[31941]=17118;
squeal_samples[31942]=13588;
squeal_samples[31943]=10276;
squeal_samples[31944]=7187;
squeal_samples[31945]=4473;
squeal_samples[31946]=5854;
squeal_samples[31947]=8770;
squeal_samples[31948]=11561;
squeal_samples[31949]=14231;
squeal_samples[31950]=16774;
squeal_samples[31951]=19222;
squeal_samples[31952]=21539;
squeal_samples[31953]=23779;
squeal_samples[31954]=25896;
squeal_samples[31955]=27942;
squeal_samples[31956]=29875;
squeal_samples[31957]=31737;
squeal_samples[31958]=33510;
squeal_samples[31959]=35201;
squeal_samples[31960]=36827;
squeal_samples[31961]=38368;
squeal_samples[31962]=39850;
squeal_samples[31963]=41254;
squeal_samples[31964]=42606;
squeal_samples[31965]=43888;
squeal_samples[31966]=45115;
squeal_samples[31967]=46290;
squeal_samples[31968]=47403;
squeal_samples[31969]=48483;
squeal_samples[31970]=49500;
squeal_samples[31971]=50474;
squeal_samples[31972]=51410;
squeal_samples[31973]=52299;
squeal_samples[31974]=53150;
squeal_samples[31975]=53960;
squeal_samples[31976]=54261;
squeal_samples[31977]=49629;
squeal_samples[31978]=44012;
squeal_samples[31979]=38754;
squeal_samples[31980]=33831;
squeal_samples[31981]=29232;
squeal_samples[31982]=24913;
squeal_samples[31983]=20880;
squeal_samples[31984]=17108;
squeal_samples[31985]=13573;
squeal_samples[31986]=10267;
squeal_samples[31987]=7173;
squeal_samples[31988]=4461;
squeal_samples[31989]=5844;
squeal_samples[31990]=8756;
squeal_samples[31991]=11550;
squeal_samples[31992]=14218;
squeal_samples[31993]=16763;
squeal_samples[31994]=19209;
squeal_samples[31995]=21530;
squeal_samples[31996]=23762;
squeal_samples[31997]=25889;
squeal_samples[31998]=27925;
squeal_samples[31999]=29867;
squeal_samples[32000]=31724;
squeal_samples[32001]=33498;
squeal_samples[32002]=35189;
squeal_samples[32003]=36814;
squeal_samples[32004]=38357;
squeal_samples[32005]=39837;
squeal_samples[32006]=41245;
squeal_samples[32007]=42591;
squeal_samples[32008]=43878;
squeal_samples[32009]=45101;
squeal_samples[32010]=46279;
squeal_samples[32011]=47391;
squeal_samples[32012]=48471;
squeal_samples[32013]=49488;
squeal_samples[32014]=50463;
squeal_samples[32015]=51396;
squeal_samples[32016]=52289;
squeal_samples[32017]=53136;
squeal_samples[32018]=53951;
squeal_samples[32019]=54246;
squeal_samples[32020]=49619;
squeal_samples[32021]=43999;
squeal_samples[32022]=38742;
squeal_samples[32023]=33820;
squeal_samples[32024]=29219;
squeal_samples[32025]=24901;
squeal_samples[32026]=20870;
squeal_samples[32027]=17093;
squeal_samples[32028]=13565;
squeal_samples[32029]=10252;
squeal_samples[32030]=7161;
squeal_samples[32031]=4453;
squeal_samples[32032]=5826;
squeal_samples[32033]=8751;
squeal_samples[32034]=11534;
squeal_samples[32035]=14207;
squeal_samples[32036]=16751;
squeal_samples[32037]=19197;
squeal_samples[32038]=21518;
squeal_samples[32039]=23750;
squeal_samples[32040]=25878;
squeal_samples[32041]=27912;
squeal_samples[32042]=29855;
squeal_samples[32043]=31713;
squeal_samples[32044]=33483;
squeal_samples[32045]=35181;
squeal_samples[32046]=36799;
squeal_samples[32047]=38348;
squeal_samples[32048]=39823;
squeal_samples[32049]=41234;
squeal_samples[32050]=42578;
squeal_samples[32051]=43866;
squeal_samples[32052]=45092;
squeal_samples[32053]=46263;
squeal_samples[32054]=47383;
squeal_samples[32055]=48457;
squeal_samples[32056]=49476;
squeal_samples[32057]=50452;
squeal_samples[32058]=51382;
squeal_samples[32059]=52279;
squeal_samples[32060]=53124;
squeal_samples[32061]=53938;
squeal_samples[32062]=54236;
squeal_samples[32063]=49604;
squeal_samples[32064]=43989;
squeal_samples[32065]=38729;
squeal_samples[32066]=33810;
squeal_samples[32067]=29204;
squeal_samples[32068]=24893;
squeal_samples[32069]=20854;
squeal_samples[32070]=17084;
squeal_samples[32071]=13551;
squeal_samples[32072]=10240;
squeal_samples[32073]=7152;
squeal_samples[32074]=4436;
squeal_samples[32075]=5819;
squeal_samples[32076]=8735;
squeal_samples[32077]=11524;
squeal_samples[32078]=14196;
squeal_samples[32079]=16737;
squeal_samples[32080]=19185;
squeal_samples[32081]=21508;
squeal_samples[32082]=23736;
squeal_samples[32083]=25868;
squeal_samples[32084]=27899;
squeal_samples[32085]=29844;
squeal_samples[32086]=31699;
squeal_samples[32087]=33474;
squeal_samples[32088]=35166;
squeal_samples[32089]=36789;
squeal_samples[32090]=38336;
squeal_samples[32091]=39809;
squeal_samples[32092]=41224;
squeal_samples[32093]=42566;
squeal_samples[32094]=43853;
squeal_samples[32095]=45080;
squeal_samples[32096]=46251;
squeal_samples[32097]=47371;
squeal_samples[32098]=48444;
squeal_samples[32099]=49467;
squeal_samples[32100]=50436;
squeal_samples[32101]=51374;
squeal_samples[32102]=52263;
squeal_samples[32103]=53114;
squeal_samples[32104]=53925;
squeal_samples[32105]=54224;
squeal_samples[32106]=49593;
squeal_samples[32107]=43977;
squeal_samples[32108]=38715;
squeal_samples[32109]=33799;
squeal_samples[32110]=29191;
squeal_samples[32111]=24882;
squeal_samples[32112]=20840;
squeal_samples[32113]=17073;
squeal_samples[32114]=13538;
squeal_samples[32115]=10227;
squeal_samples[32116]=7141;
squeal_samples[32117]=4649;
squeal_samples[32118]=6516;
squeal_samples[32119]=9393;
squeal_samples[32120]=12156;
squeal_samples[32121]=14793;
squeal_samples[32122]=17321;
squeal_samples[32123]=19731;
squeal_samples[32124]=22030;
squeal_samples[32125]=24238;
squeal_samples[32126]=26346;
squeal_samples[32127]=28356;
squeal_samples[32128]=30281;
squeal_samples[32129]=32117;
squeal_samples[32130]=33872;
squeal_samples[32131]=35552;
squeal_samples[32132]=37150;
squeal_samples[32133]=38677;
squeal_samples[32134]=40134;
squeal_samples[32135]=41537;
squeal_samples[32136]=42862;
squeal_samples[32137]=44136;
squeal_samples[32138]=45349;
squeal_samples[32139]=46511;
squeal_samples[32140]=47619;
squeal_samples[32141]=48677;
squeal_samples[32142]=49686;
squeal_samples[32143]=50656;
squeal_samples[32144]=51570;
squeal_samples[32145]=52455;
squeal_samples[32146]=53296;
squeal_samples[32147]=54105;
squeal_samples[32148]=54021;
squeal_samples[32149]=48935;
squeal_samples[32150]=43361;
squeal_samples[32151]=38139;
squeal_samples[32152]=33261;
squeal_samples[32153]=28684;
squeal_samples[32154]=24403;
squeal_samples[32155]=20401;
squeal_samples[32156]=16653;
squeal_samples[32157]=13145;
squeal_samples[32158]=9866;
squeal_samples[32159]=6792;
squeal_samples[32160]=4335;
squeal_samples[32161]=6199;
squeal_samples[32162]=9105;
squeal_samples[32163]=11868;
squeal_samples[32164]=14524;
squeal_samples[32165]=17058;
squeal_samples[32166]=19484;
squeal_samples[32167]=21800;
squeal_samples[32168]=24011;
squeal_samples[32169]=26124;
squeal_samples[32170]=28149;
squeal_samples[32171]=30078;
squeal_samples[32172]=31927;
squeal_samples[32173]=33687;
squeal_samples[32174]=35371;
squeal_samples[32175]=36982;
squeal_samples[32176]=38518;
squeal_samples[32177]=39981;
squeal_samples[32178]=41384;
squeal_samples[32179]=42720;
squeal_samples[32180]=43999;
squeal_samples[32181]=45218;
squeal_samples[32182]=46386;
squeal_samples[32183]=47497;
squeal_samples[32184]=48563;
squeal_samples[32185]=49576;
squeal_samples[32186]=50546;
squeal_samples[32187]=51472;
squeal_samples[32188]=52361;
squeal_samples[32189]=53203;
squeal_samples[32190]=54011;
squeal_samples[32191]=53935;
squeal_samples[32192]=48849;
squeal_samples[32193]=43287;
squeal_samples[32194]=38066;
squeal_samples[32195]=33189;
squeal_samples[32196]=28618;
squeal_samples[32197]=24343;
squeal_samples[32198]=20337;
squeal_samples[32199]=16601;
squeal_samples[32200]=13092;
squeal_samples[32201]=9816;
squeal_samples[32202]=6744;
squeal_samples[32203]=4595;
squeal_samples[32204]=6861;
squeal_samples[32205]=9728;
squeal_samples[32206]=12473;
squeal_samples[32207]=15097;
squeal_samples[32208]=17605;
squeal_samples[32209]=20000;
squeal_samples[32210]=22296;
squeal_samples[32211]=24483;
squeal_samples[32212]=26579;
squeal_samples[32213]=28581;
squeal_samples[32214]=30491;
squeal_samples[32215]=32319;
squeal_samples[32216]=34063;
squeal_samples[32217]=35731;
squeal_samples[32218]=37325;
squeal_samples[32219]=38840;
squeal_samples[32220]=40296;
squeal_samples[32221]=41680;
squeal_samples[32222]=43002;
squeal_samples[32223]=44269;
squeal_samples[32224]=45478;
squeal_samples[32225]=46628;
squeal_samples[32226]=47729;
squeal_samples[32227]=48786;
squeal_samples[32228]=49785;
squeal_samples[32229]=50753;
squeal_samples[32230]=51660;
squeal_samples[32231]=52540;
squeal_samples[32232]=53374;
squeal_samples[32233]=54183;
squeal_samples[32234]=53613;
squeal_samples[32235]=48203;
squeal_samples[32236]=42666;
squeal_samples[32237]=37492;
squeal_samples[32238]=32649;
squeal_samples[32239]=28109;
squeal_samples[32240]=23867;
squeal_samples[32241]=19894;
squeal_samples[32242]=16178;
squeal_samples[32243]=12704;
squeal_samples[32244]=9450;
squeal_samples[32245]=6401;
squeal_samples[32246]=4274;
squeal_samples[32247]=6550;
squeal_samples[32248]=9429;
squeal_samples[32249]=12192;
squeal_samples[32250]=14822;
squeal_samples[32251]=17345;
squeal_samples[32252]=19754;
squeal_samples[32253]=22056;
squeal_samples[32254]=24256;
squeal_samples[32255]=26358;
squeal_samples[32256]=28371;
squeal_samples[32257]=30287;
squeal_samples[32258]=32125;
squeal_samples[32259]=33875;
squeal_samples[32260]=35553;
squeal_samples[32261]=37153;
squeal_samples[32262]=38679;
squeal_samples[32263]=40135;
squeal_samples[32264]=41536;
squeal_samples[32265]=42856;
squeal_samples[32266]=44136;
squeal_samples[32267]=45342;
squeal_samples[32268]=46505;
squeal_samples[32269]=47609;
squeal_samples[32270]=48668;
squeal_samples[32271]=49679;
squeal_samples[32272]=50639;
squeal_samples[32273]=51564;
squeal_samples[32274]=52439;
squeal_samples[32275]=53283;
squeal_samples[32276]=54083;
squeal_samples[32277]=54005;
squeal_samples[32278]=48917;
squeal_samples[32279]=43345;
squeal_samples[32280]=38117;
squeal_samples[32281]=33237;
squeal_samples[32282]=28658;
squeal_samples[32283]=24384;
squeal_samples[32284]=20376;
squeal_samples[32285]=16626;
squeal_samples[32286]=13124;
squeal_samples[32287]=9836;
squeal_samples[32288]=6772;
squeal_samples[32289]=4299;
squeal_samples[32290]=6180;
squeal_samples[32291]=9072;
squeal_samples[32292]=11851;
squeal_samples[32293]=14493;
squeal_samples[32294]=17037;
squeal_samples[32295]=19451;
squeal_samples[32296]=21770;
squeal_samples[32297]=23981;
squeal_samples[32298]=26093;
squeal_samples[32299]=28119;
squeal_samples[32300]=30047;
squeal_samples[32301]=31897;
squeal_samples[32302]=33656;
squeal_samples[32303]=35340;
squeal_samples[32304]=36947;
squeal_samples[32305]=38481;
squeal_samples[32306]=39952;
squeal_samples[32307]=41351;
squeal_samples[32308]=42692;
squeal_samples[32309]=43967;
squeal_samples[32310]=45188;
squeal_samples[32311]=46355;
squeal_samples[32312]=47466;
squeal_samples[32313]=48528;
squeal_samples[32314]=49540;
squeal_samples[32315]=50514;
squeal_samples[32316]=51438;
squeal_samples[32317]=52322;
squeal_samples[32318]=53169;
squeal_samples[32319]=53979;
squeal_samples[32320]=54271;
squeal_samples[32321]=49634;
squeal_samples[32322]=44005;
squeal_samples[32323]=38747;
squeal_samples[32324]=33816;
squeal_samples[32325]=29211;
squeal_samples[32326]=24888;
squeal_samples[32327]=20856;
squeal_samples[32328]=17070;
squeal_samples[32329]=13538;
squeal_samples[32330]=10230;
squeal_samples[32331]=7131;
squeal_samples[32332]=4415;
squeal_samples[32333]=5795;
squeal_samples[32334]=8707;
squeal_samples[32335]=11489;
squeal_samples[32336]=14162;
squeal_samples[32337]=16705;
squeal_samples[32338]=19144;
squeal_samples[32339]=21473;
squeal_samples[32340]=23699;
squeal_samples[32341]=25825;
squeal_samples[32342]=27858;
squeal_samples[32343]=29797;
squeal_samples[32344]=31654;
squeal_samples[32345]=33430;
squeal_samples[32346]=35120;
squeal_samples[32347]=36740;
squeal_samples[32348]=38284;
squeal_samples[32349]=39761;
squeal_samples[32350]=41165;
squeal_samples[32351]=42513;
squeal_samples[32352]=43796;
squeal_samples[32353]=45025;
squeal_samples[32354]=46195;
squeal_samples[32355]=47320;
squeal_samples[32356]=48383;
squeal_samples[32357]=49406;
squeal_samples[32358]=50381;
squeal_samples[32359]=51311;
squeal_samples[32360]=52203;
squeal_samples[32361]=53051;
squeal_samples[32362]=53870;
squeal_samples[32363]=54434;
squeal_samples[32364]=50347;
squeal_samples[32365]=44680;
squeal_samples[32366]=39373;
squeal_samples[32367]=34404;
squeal_samples[32368]=29756;
squeal_samples[32369]=25401;
squeal_samples[32370]=21328;
squeal_samples[32371]=17521;
squeal_samples[32372]=13957;
squeal_samples[32373]=10616;
squeal_samples[32374]=7499;
squeal_samples[32375]=4616;
squeal_samples[32376]=5410;
squeal_samples[32377]=8339;
squeal_samples[32378]=11139;
squeal_samples[32379]=13819;
squeal_samples[32380]=16388;
squeal_samples[32381]=18829;
squeal_samples[32382]=21176;
squeal_samples[32383]=23413;
squeal_samples[32384]=25555;
squeal_samples[32385]=27600;
squeal_samples[32386]=29550;
squeal_samples[32387]=31417;
squeal_samples[32388]=33197;
squeal_samples[32389]=34906;
squeal_samples[32390]=36529;
squeal_samples[32391]=38083;
squeal_samples[32392]=39565;
squeal_samples[32393]=40984;
squeal_samples[32394]=42338;
squeal_samples[32395]=43626;
squeal_samples[32396]=44866;
squeal_samples[32397]=46044;
squeal_samples[32398]=47164;
squeal_samples[32399]=48243;
squeal_samples[32400]=49265;
squeal_samples[32401]=50252;
squeal_samples[32402]=51184;
squeal_samples[32403]=52082;
squeal_samples[32404]=52935;
squeal_samples[32405]=53754;
squeal_samples[32406]=54485;
squeal_samples[32407]=51076;
squeal_samples[32408]=45356;
squeal_samples[32409]=40008;
squeal_samples[32410]=34994;
squeal_samples[32411]=30308;
squeal_samples[32412]=25920;
squeal_samples[32413]=21811;
squeal_samples[32414]=17970;
squeal_samples[32415]=14377;
squeal_samples[32416]=11008;
squeal_samples[32417]=7863;
squeal_samples[32418]=4960;
squeal_samples[32419]=5732;
squeal_samples[32420]=8647;
squeal_samples[32421]=11436;
squeal_samples[32422]=14100;
squeal_samples[32423]=16656;
squeal_samples[32424]=19092;
squeal_samples[32425]=21414;
squeal_samples[32426]=23650;
squeal_samples[32427]=25770;
squeal_samples[32428]=27813;
squeal_samples[32429]=29750;
squeal_samples[32430]=31611;
squeal_samples[32431]=33380;
squeal_samples[32432]=35077;
squeal_samples[32433]=36696;
squeal_samples[32434]=38239;
squeal_samples[32435]=39716;
squeal_samples[32436]=41123;
squeal_samples[32437]=42473;
squeal_samples[32438]=43755;
squeal_samples[32439]=44989;
squeal_samples[32440]=46161;
squeal_samples[32441]=47278;
squeal_samples[32442]=48349;
squeal_samples[32443]=49369;
squeal_samples[32444]=50347;
squeal_samples[32445]=51275;
squeal_samples[32446]=52168;
squeal_samples[32447]=53021;
squeal_samples[32448]=53834;
squeal_samples[32449]=54399;
squeal_samples[32450]=50317;
squeal_samples[32451]=44646;
squeal_samples[32452]=39335;
squeal_samples[32453]=34377;
squeal_samples[32454]=29723;
squeal_samples[32455]=25372;
squeal_samples[32456]=21299;
squeal_samples[32457]=17490;
squeal_samples[32458]=13926;
squeal_samples[32459]=10587;
squeal_samples[32460]=7467;
squeal_samples[32461]=4722;
squeal_samples[32462]=6088;
squeal_samples[32463]=8985;
squeal_samples[32464]=11762;
squeal_samples[32465]=14408;
squeal_samples[32466]=16947;
squeal_samples[32467]=19374;
squeal_samples[32468]=21685;
squeal_samples[32469]=23901;
squeal_samples[32470]=26018;
squeal_samples[32471]=28039;
squeal_samples[32472]=29977;
squeal_samples[32473]=31821;
squeal_samples[32474]=33589;
squeal_samples[32475]=35269;
squeal_samples[32476]=36881;
squeal_samples[32477]=38416;
squeal_samples[32478]=39882;
squeal_samples[32479]=41285;
squeal_samples[32480]=42624;
squeal_samples[32481]=43898;
squeal_samples[32482]=45128;
squeal_samples[32483]=46284;
squeal_samples[32484]=47407;
squeal_samples[32485]=48463;
squeal_samples[32486]=49484;
squeal_samples[32487]=50452;
squeal_samples[32488]=51379;
squeal_samples[32489]=52263;
squeal_samples[32490]=53107;
squeal_samples[32491]=53921;
squeal_samples[32492]=54476;
squeal_samples[32493]=50394;
squeal_samples[32494]=44718;
squeal_samples[32495]=39408;
squeal_samples[32496]=34432;
squeal_samples[32497]=29778;
squeal_samples[32498]=25425;
squeal_samples[32499]=21344;
squeal_samples[32500]=17537;
squeal_samples[32501]=13964;
squeal_samples[32502]=10627;
squeal_samples[32503]=7497;
squeal_samples[32504]=4620;
squeal_samples[32505]=5411;
squeal_samples[32506]=8334;
squeal_samples[32507]=11134;
squeal_samples[32508]=13818;
squeal_samples[32509]=16379;
squeal_samples[32510]=18831;
squeal_samples[32511]=21162;
squeal_samples[32512]=23400;
squeal_samples[32513]=25540;
squeal_samples[32514]=27582;
squeal_samples[32515]=29540;
squeal_samples[32516]=31403;
squeal_samples[32517]=33186;
squeal_samples[32518]=34887;
squeal_samples[32519]=36512;
squeal_samples[32520]=38061;
squeal_samples[32521]=39550;
squeal_samples[32522]=40964;
squeal_samples[32523]=42317;
squeal_samples[32524]=43606;
squeal_samples[32525]=44841;
squeal_samples[32526]=46015;
squeal_samples[32527]=47148;
squeal_samples[32528]=48218;
squeal_samples[32529]=49249;
squeal_samples[32530]=50221;
squeal_samples[32531]=51168;
squeal_samples[32532]=52051;
squeal_samples[32533]=52916;
squeal_samples[32534]=53720;
squeal_samples[32535]=54514;
squeal_samples[32536]=51871;
squeal_samples[32537]=46105;
squeal_samples[32538]=40704;
squeal_samples[32539]=35645;
squeal_samples[32540]=30920;
squeal_samples[32541]=26485;
squeal_samples[32542]=22340;
squeal_samples[32543]=18465;
squeal_samples[32544]=14835;
squeal_samples[32545]=11433;
squeal_samples[32546]=8256;
squeal_samples[32547]=5283;
squeal_samples[32548]=4696;
squeal_samples[32549]=7609;
squeal_samples[32550]=10445;
squeal_samples[32551]=13150;
squeal_samples[32552]=15745;
squeal_samples[32553]=18221;
squeal_samples[32554]=20577;
squeal_samples[32555]=22851;
squeal_samples[32556]=25004;
squeal_samples[32557]=27083;
squeal_samples[32558]=29046;
squeal_samples[32559]=30937;
squeal_samples[32560]=32739;
squeal_samples[32561]=34457;
squeal_samples[32562]=36103;
squeal_samples[32563]=37675;
squeal_samples[32564]=39173;
squeal_samples[32565]=40606;
squeal_samples[32566]=41972;
squeal_samples[32567]=43282;
squeal_samples[32568]=44526;
squeal_samples[32569]=45724;
squeal_samples[32570]=46855;
squeal_samples[32571]=47949;
squeal_samples[32572]=48984;
squeal_samples[32573]=49972;
squeal_samples[32574]=50925;
squeal_samples[32575]=51824;
squeal_samples[32576]=52692;
squeal_samples[32577]=53517;
squeal_samples[32578]=54311;
squeal_samples[32579]=53149;
squeal_samples[32580]=47505;
squeal_samples[32581]=42010;
squeal_samples[32582]=36868;
squeal_samples[32583]=32057;
squeal_samples[32584]=27553;
squeal_samples[32585]=23343;
squeal_samples[32586]=19397;
squeal_samples[32587]=15709;
squeal_samples[32588]=12250;
squeal_samples[32589]=9023;
squeal_samples[32590]=5997;
squeal_samples[32591]=4292;
squeal_samples[32592]=6870;
squeal_samples[32593]=9733;
squeal_samples[32594]=12475;
squeal_samples[32595]=15093;
squeal_samples[32596]=17602;
squeal_samples[32597]=19985;
squeal_samples[32598]=22281;
squeal_samples[32599]=24465;
squeal_samples[32600]=26556;
squeal_samples[32601]=28553;
squeal_samples[32602]=30462;
squeal_samples[32603]=32288;
squeal_samples[32604]=34026;
squeal_samples[32605]=35690;
squeal_samples[32606]=37275;
squeal_samples[32607]=38795;
squeal_samples[32608]=40238;
squeal_samples[32609]=41631;
squeal_samples[32610]=42947;
squeal_samples[32611]=44211;
squeal_samples[32612]=45419;
squeal_samples[32613]=46565;
squeal_samples[32614]=47666;
squeal_samples[32615]=48715;
squeal_samples[32616]=49722;
squeal_samples[32617]=50678;
squeal_samples[32618]=51590;
squeal_samples[32619]=52466;
squeal_samples[32620]=53299;
squeal_samples[32621]=54099;
squeal_samples[32622]=54015;
squeal_samples[32623]=48918;
squeal_samples[32624]=43337;
squeal_samples[32625]=38108;
squeal_samples[32626]=33224;
squeal_samples[32627]=28637;
squeal_samples[32628]=24357;
squeal_samples[32629]=20341;
squeal_samples[32630]=16596;
squeal_samples[32631]=13083;
squeal_samples[32632]=9794;
squeal_samples[32633]=6722;
squeal_samples[32634]=4251;
squeal_samples[32635]=6123;
squeal_samples[32636]=9021;
squeal_samples[32637]=11787;
squeal_samples[32638]=14436;
squeal_samples[32639]=16974;
squeal_samples[32640]=19394;
squeal_samples[32641]=21702;
squeal_samples[32642]=23917;
squeal_samples[32643]=26026;
squeal_samples[32644]=28054;
squeal_samples[32645]=29976;
squeal_samples[32646]=31826;
squeal_samples[32647]=33584;
squeal_samples[32648]=35271;
squeal_samples[32649]=36873;
squeal_samples[32650]=38411;
squeal_samples[32651]=39876;
squeal_samples[32652]=41273;
squeal_samples[32653]=42612;
squeal_samples[32654]=43888;
squeal_samples[32655]=45107;
squeal_samples[32656]=46273;
squeal_samples[32657]=47384;
squeal_samples[32658]=48445;
squeal_samples[32659]=49458;
squeal_samples[32660]=50433;
squeal_samples[32661]=51353;
squeal_samples[32662]=52237;
squeal_samples[32663]=53085;
squeal_samples[32664]=53890;
squeal_samples[32665]=54453;
squeal_samples[32666]=50361;
squeal_samples[32667]=44688;
squeal_samples[32668]=39373;
squeal_samples[32669]=34400;
squeal_samples[32670]=29744;
squeal_samples[32671]=25385;
squeal_samples[32672]=21307;
squeal_samples[32673]=17496;
squeal_samples[32674]=13927;
squeal_samples[32675]=10588;
squeal_samples[32676]=7456;
squeal_samples[32677]=4584;
squeal_samples[32678]=5363;
squeal_samples[32679]=8298;
squeal_samples[32680]=11093;
squeal_samples[32681]=13775;
squeal_samples[32682]=16334;
squeal_samples[32683]=18786;
squeal_samples[32684]=21119;
squeal_samples[32685]=23360;
squeal_samples[32686]=25501;
squeal_samples[32687]=27538;
squeal_samples[32688]=29496;
squeal_samples[32689]=31358;
squeal_samples[32690]=33142;
squeal_samples[32691]=34843;
squeal_samples[32692]=36465;
squeal_samples[32693]=38020;
squeal_samples[32694]=39502;
squeal_samples[32695]=40917;
squeal_samples[32696]=42271;
squeal_samples[32697]=43562;
squeal_samples[32698]=44797;
squeal_samples[32699]=45969;
squeal_samples[32700]=47098;
squeal_samples[32701]=48170;
squeal_samples[32702]=49196;
squeal_samples[32703]=50181;
squeal_samples[32704]=51113;
squeal_samples[32705]=52011;
squeal_samples[32706]=52866;
squeal_samples[32707]=53681;
squeal_samples[32708]=54466;
squeal_samples[32709]=51826;
squeal_samples[32710]=46063;
squeal_samples[32711]=40649;
squeal_samples[32712]=35601;
squeal_samples[32713]=30865;
squeal_samples[32714]=26437;
squeal_samples[32715]=22288;
squeal_samples[32716]=18416;
squeal_samples[32717]=14784;
squeal_samples[32718]=11388;
squeal_samples[32719]=8206;
squeal_samples[32720]=5231;
squeal_samples[32721]=5321;
squeal_samples[32722]=8242;
squeal_samples[32723]=11052;
squeal_samples[32724]=13724;
squeal_samples[32725]=16294;
squeal_samples[32726]=18742;
squeal_samples[32727]=21080;
squeal_samples[32728]=23322;
squeal_samples[32729]=25457;
squeal_samples[32730]=27509;
squeal_samples[32731]=29455;
squeal_samples[32732]=31329;
squeal_samples[32733]=33104;
squeal_samples[32734]=34811;
squeal_samples[32735]=36435;
squeal_samples[32736]=37991;
squeal_samples[32737]=39467;
squeal_samples[32738]=40889;
squeal_samples[32739]=42241;
squeal_samples[32740]=43534;
squeal_samples[32741]=44767;
squeal_samples[32742]=45947;
squeal_samples[32743]=47074;
squeal_samples[32744]=48145;
squeal_samples[32745]=49175;
squeal_samples[32746]=50155;
squeal_samples[32747]=51091;
squeal_samples[32748]=51988;
squeal_samples[32749]=52841;
squeal_samples[32750]=53659;
squeal_samples[32751]=54440;
squeal_samples[32752]=51806;
squeal_samples[32753]=46036;
squeal_samples[32754]=40634;
squeal_samples[32755]=35581;
squeal_samples[32756]=30847;
squeal_samples[32757]=26420;
squeal_samples[32758]=22268;
squeal_samples[32759]=18400;
squeal_samples[32760]=14765;
squeal_samples[32761]=11370;
squeal_samples[32762]=8194;
squeal_samples[32763]=5217;
squeal_samples[32764]=5302;
squeal_samples[32765]=8233;
squeal_samples[32766]=11030;
squeal_samples[32767]=13715;
squeal_samples[32768]=16278;
squeal_samples[32769]=18725;
squeal_samples[32770]=21069;
squeal_samples[32771]=23301;
squeal_samples[32772]=25448;
squeal_samples[32773]=27488;
squeal_samples[32774]=29439;
squeal_samples[32775]=31311;
squeal_samples[32776]=33089;
squeal_samples[32777]=34796;
squeal_samples[32778]=36416;
squeal_samples[32779]=37972;
squeal_samples[32780]=39457;
squeal_samples[32781]=40873;
squeal_samples[32782]=42226;
squeal_samples[32783]=43521;
squeal_samples[32784]=44752;
squeal_samples[32785]=45932;
squeal_samples[32786]=47058;
squeal_samples[32787]=48136;
squeal_samples[32788]=49160;
squeal_samples[32789]=50139;
squeal_samples[32790]=51076;
squeal_samples[32791]=51972;
squeal_samples[32792]=52826;
squeal_samples[32793]=53649;
squeal_samples[32794]=54425;
squeal_samples[32795]=51796;
squeal_samples[32796]=46022;
squeal_samples[32797]=40622;
squeal_samples[32798]=35567;
squeal_samples[32799]=30836;
squeal_samples[32800]=26405;
squeal_samples[32801]=22260;
squeal_samples[32802]=18382;
squeal_samples[32803]=14756;
squeal_samples[32804]=11356;
squeal_samples[32805]=8180;
squeal_samples[32806]=5202;
squeal_samples[32807]=5288;
squeal_samples[32808]=8219;
squeal_samples[32809]=11020;
squeal_samples[32810]=13699;
squeal_samples[32811]=16269;
squeal_samples[32812]=18711;
squeal_samples[32813]=21056;
squeal_samples[32814]=23288;
squeal_samples[32815]=25431;
squeal_samples[32816]=27472;
squeal_samples[32817]=29432;
squeal_samples[32818]=31292;
squeal_samples[32819]=33083;
squeal_samples[32820]=34777;
squeal_samples[32821]=36406;
squeal_samples[32822]=37958;
squeal_samples[32823]=39446;
squeal_samples[32824]=40859;
squeal_samples[32825]=42215;
squeal_samples[32826]=43505;
squeal_samples[32827]=44743;
squeal_samples[32828]=45916;
squeal_samples[32829]=47048;
squeal_samples[32830]=48121;
squeal_samples[32831]=49149;
squeal_samples[32832]=50123;
squeal_samples[32833]=51068;
squeal_samples[32834]=51954;
squeal_samples[32835]=52817;
squeal_samples[32836]=53633;
squeal_samples[32837]=54414;
squeal_samples[32838]=52564;
squeal_samples[32839]=46798;
squeal_samples[32840]=41342;
squeal_samples[32841]=36245;
squeal_samples[32842]=31464;
squeal_samples[32843]=26996;
squeal_samples[32844]=22809;
squeal_samples[32845]=18901;
squeal_samples[32846]=15233;
squeal_samples[32847]=11809;
squeal_samples[32848]=8596;
squeal_samples[32849]=5597;
squeal_samples[32850]=4407;
squeal_samples[32851]=7196;
squeal_samples[32852]=10044;
squeal_samples[32853]=12766;
squeal_samples[32854]=15368;
squeal_samples[32855]=17860;
squeal_samples[32856]=20233;
squeal_samples[32857]=22506;
squeal_samples[32858]=24685;
squeal_samples[32859]=26755;
squeal_samples[32860]=28743;
squeal_samples[32861]=30644;
squeal_samples[32862]=32446;
squeal_samples[32863]=34184;
squeal_samples[32864]=35831;
squeal_samples[32865]=37416;
squeal_samples[32866]=38921;
squeal_samples[32867]=40361;
squeal_samples[32868]=41736;
squeal_samples[32869]=43053;
squeal_samples[32870]=44302;
squeal_samples[32871]=45500;
squeal_samples[32872]=46643;
squeal_samples[32873]=47740;
squeal_samples[32874]=48781;
squeal_samples[32875]=49777;
squeal_samples[32876]=50725;
squeal_samples[32877]=51639;
squeal_samples[32878]=52507;
squeal_samples[32879]=53333;
squeal_samples[32880]=54136;
squeal_samples[32881]=54033;
squeal_samples[32882]=48942;
squeal_samples[32883]=43351;
squeal_samples[32884]=38122;
squeal_samples[32885]=33221;
squeal_samples[32886]=28639;
squeal_samples[32887]=24351;
squeal_samples[32888]=20330;
squeal_samples[32889]=16579;
squeal_samples[32890]=13062;
squeal_samples[32891]=9771;
squeal_samples[32892]=6696;
squeal_samples[32893]=4223;
squeal_samples[32894]=6090;
squeal_samples[32895]=8984;
squeal_samples[32896]=11753;
squeal_samples[32897]=14399;
squeal_samples[32898]=16929;
squeal_samples[32899]=19352;
squeal_samples[32900]=21657;
squeal_samples[32901]=23874;
squeal_samples[32902]=25983;
squeal_samples[32903]=28003;
squeal_samples[32904]=29929;
squeal_samples[32905]=31776;
squeal_samples[32906]=33530;
squeal_samples[32907]=35216;
squeal_samples[32908]=36819;
squeal_samples[32909]=38357;
squeal_samples[32910]=39819;
squeal_samples[32911]=41222;
squeal_samples[32912]=42554;
squeal_samples[32913]=43831;
squeal_samples[32914]=45051;
squeal_samples[32915]=46212;
squeal_samples[32916]=47325;
squeal_samples[32917]=48384;
squeal_samples[32918]=49399;
squeal_samples[32919]=50366;
squeal_samples[32920]=51288;
squeal_samples[32921]=52177;
squeal_samples[32922]=53018;
squeal_samples[32923]=53826;
squeal_samples[32924]=54547;
squeal_samples[32925]=51119;
squeal_samples[32926]=45392;
squeal_samples[32927]=40031;
squeal_samples[32928]=35007;
squeal_samples[32929]=30308;
squeal_samples[32930]=25913;
squeal_samples[32931]=21794;
squeal_samples[32932]=17947;
squeal_samples[32933]=14339;
squeal_samples[32934]=10967;
squeal_samples[32935]=7811;
squeal_samples[32936]=4858;
squeal_samples[32937]=4963;
squeal_samples[32938]=7904;
squeal_samples[32939]=10714;
squeal_samples[32940]=13410;
squeal_samples[32941]=15980;
squeal_samples[32942]=18445;
squeal_samples[32943]=20790;
squeal_samples[32944]=23044;
squeal_samples[32945]=25185;
squeal_samples[32946]=27251;
squeal_samples[32947]=29203;
squeal_samples[32948]=31083;
squeal_samples[32949]=32876;
squeal_samples[32950]=34579;
squeal_samples[32951]=36219;
squeal_samples[32952]=37772;
squeal_samples[32953]=39265;
squeal_samples[32954]=40688;
squeal_samples[32955]=42046;
squeal_samples[32956]=43348;
squeal_samples[32957]=44586;
squeal_samples[32958]=45771;
squeal_samples[32959]=46902;
squeal_samples[32960]=47976;
squeal_samples[32961]=49016;
squeal_samples[32962]=49990;
squeal_samples[32963]=50937;
squeal_samples[32964]=51835;
squeal_samples[32965]=52696;
squeal_samples[32966]=53512;
squeal_samples[32967]=54299;
squeal_samples[32968]=53140;
squeal_samples[32969]=47480;
squeal_samples[32970]=41985;
squeal_samples[32971]=36839;
squeal_samples[32972]=32024;
squeal_samples[32973]=27516;
squeal_samples[32974]=23292;
squeal_samples[32975]=19350;
squeal_samples[32976]=15652;
squeal_samples[32977]=12193;
squeal_samples[32978]=8959;
squeal_samples[32979]=5934;
squeal_samples[32980]=4226;
squeal_samples[32981]=6804;
squeal_samples[32982]=9663;
squeal_samples[32983]=12403;
squeal_samples[32984]=15016;
squeal_samples[32985]=17527;
squeal_samples[32986]=19908;
squeal_samples[32987]=22198;
squeal_samples[32988]=24385;
squeal_samples[32989]=26471;
squeal_samples[32990]=28474;
squeal_samples[32991]=30373;
squeal_samples[32992]=32200;
squeal_samples[32993]=33934;
squeal_samples[32994]=35602;
squeal_samples[32995]=37184;
squeal_samples[32996]=38704;
squeal_samples[32997]=40147;
squeal_samples[32998]=41532;
squeal_samples[32999]=42853;
squeal_samples[33000]=44116;
squeal_samples[33001]=45316;
squeal_samples[33002]=46469;
squeal_samples[33003]=47566;
squeal_samples[33004]=48617;
squeal_samples[33005]=49619;
squeal_samples[33006]=50571;
squeal_samples[33007]=51494;
squeal_samples[33008]=52358;
squeal_samples[33009]=53203;
squeal_samples[33010]=53995;
squeal_samples[33011]=54277;
squeal_samples[33012]=49626;
squeal_samples[33013]=43991;
squeal_samples[33014]=38716;
squeal_samples[33015]=33783;
squeal_samples[33016]=29157;
squeal_samples[33017]=24833;
squeal_samples[33018]=20780;
squeal_samples[33019]=16996;
squeal_samples[33020]=13450;
squeal_samples[33021]=10138;
squeal_samples[33022]=7026;
squeal_samples[33023]=4535;
squeal_samples[33024]=6386;
squeal_samples[33025]=9264;
squeal_samples[33026]=12020;
squeal_samples[33027]=14651;
squeal_samples[33028]=17174;
squeal_samples[33029]=19583;
squeal_samples[33030]=21879;
squeal_samples[33031]=24078;
squeal_samples[33032]=26179;
squeal_samples[33033]=28185;
squeal_samples[33034]=30108;
squeal_samples[33035]=31942;
squeal_samples[33036]=33687;
squeal_samples[33037]=35362;
squeal_samples[33038]=36958;
squeal_samples[33039]=38486;
squeal_samples[33040]=39944;
squeal_samples[33041]=41333;
squeal_samples[33042]=42663;
squeal_samples[33043]=43933;
squeal_samples[33044]=45141;
squeal_samples[33045]=46305;
squeal_samples[33046]=47404;
squeal_samples[33047]=48465;
squeal_samples[33048]=49473;
squeal_samples[33049]=50437;
squeal_samples[33050]=51351;
squeal_samples[33051]=52237;
squeal_samples[33052]=53070;
squeal_samples[33053]=53881;
squeal_samples[33054]=54432;
squeal_samples[33055]=50335;
squeal_samples[33056]=44657;
squeal_samples[33057]=39341;
squeal_samples[33058]=34357;
squeal_samples[33059]=29703;
squeal_samples[33060]=25332;
squeal_samples[33061]=21258;
squeal_samples[33062]=17438;
squeal_samples[33063]=13867;
squeal_samples[33064]=10519;
squeal_samples[33065]=7392;
squeal_samples[33066]=4643;
squeal_samples[33067]=6002;
squeal_samples[33068]=8895;
squeal_samples[33069]=11665;
squeal_samples[33070]=14313;
squeal_samples[33071]=16851;
squeal_samples[33072]=19271;
squeal_samples[33073]=21580;
squeal_samples[33074]=23791;
squeal_samples[33075]=25908;
squeal_samples[33076]=27921;
squeal_samples[33077]=29858;
squeal_samples[33078]=31697;
squeal_samples[33079]=33462;
squeal_samples[33080]=35139;
squeal_samples[33081]=36747;
squeal_samples[33082]=38282;
squeal_samples[33083]=39746;
squeal_samples[33084]=41147;
squeal_samples[33085]=42489;
squeal_samples[33086]=43758;
squeal_samples[33087]=44987;
squeal_samples[33088]=46140;
squeal_samples[33089]=47260;
squeal_samples[33090]=48319;
squeal_samples[33091]=49337;
squeal_samples[33092]=50302;
squeal_samples[33093]=51227;
squeal_samples[33094]=52112;
squeal_samples[33095]=52956;
squeal_samples[33096]=53763;
squeal_samples[33097]=54483;
squeal_samples[33098]=51063;
squeal_samples[33099]=45329;
squeal_samples[33100]=39965;
squeal_samples[33101]=34953;
squeal_samples[33102]=30248;
squeal_samples[33103]=25856;
squeal_samples[33104]=21737;
squeal_samples[33105]=17887;
squeal_samples[33106]=14283;
squeal_samples[33107]=10910;
squeal_samples[33108]=7755;
squeal_samples[33109]=4854;
squeal_samples[33110]=5610;
squeal_samples[33111]=8533;
squeal_samples[33112]=11307;
squeal_samples[33113]=13980;
squeal_samples[33114]=16520;
squeal_samples[33115]=18960;
squeal_samples[33116]=21285;
squeal_samples[33117]=23507;
squeal_samples[33118]=25633;
squeal_samples[33119]=27665;
squeal_samples[33120]=29606;
squeal_samples[33121]=31456;
squeal_samples[33122]=33233;
squeal_samples[33123]=34918;
squeal_samples[33124]=36540;
squeal_samples[33125]=38085;
squeal_samples[33126]=39552;
squeal_samples[33127]=40969;
squeal_samples[33128]=42309;
squeal_samples[33129]=43593;
squeal_samples[33130]=44817;
squeal_samples[33131]=45990;
squeal_samples[33132]=47109;
squeal_samples[33133]=48176;
squeal_samples[33134]=49200;
squeal_samples[33135]=50169;
squeal_samples[33136]=51099;
squeal_samples[33137]=51992;
squeal_samples[33138]=52839;
squeal_samples[33139]=53651;
squeal_samples[33140]=54428;
squeal_samples[33141]=51787;
squeal_samples[33142]=46012;
squeal_samples[33143]=40606;
squeal_samples[33144]=35544;
squeal_samples[33145]=30810;
squeal_samples[33146]=26371;
squeal_samples[33147]=22226;
squeal_samples[33148]=18341;
squeal_samples[33149]=14709;
squeal_samples[33150]=11308;
squeal_samples[33151]=8127;
squeal_samples[33152]=5145;
squeal_samples[33153]=5229;
squeal_samples[33154]=8160;
squeal_samples[33155]=10957;
squeal_samples[33156]=13636;
squeal_samples[33157]=16202;
squeal_samples[33158]=18646;
squeal_samples[33159]=20985;
squeal_samples[33160]=23217;
squeal_samples[33161]=25359;
squeal_samples[33162]=27404;
squeal_samples[33163]=29357;
squeal_samples[33164]=31219;
squeal_samples[33165]=33003;
squeal_samples[33166]=34703;
squeal_samples[33167]=36330;
squeal_samples[33168]=37881;
squeal_samples[33169]=39363;
squeal_samples[33170]=40778;
squeal_samples[33171]=42132;
squeal_samples[33172]=43418;
squeal_samples[33173]=44656;
squeal_samples[33174]=45834;
squeal_samples[33175]=46959;
squeal_samples[33176]=48037;
squeal_samples[33177]=49055;
squeal_samples[33178]=50044;
squeal_samples[33179]=50967;
squeal_samples[33180]=51872;
squeal_samples[33181]=52721;
squeal_samples[33182]=53541;
squeal_samples[33183]=54318;
squeal_samples[33184]=53159;
squeal_samples[33185]=47489;
squeal_samples[33186]=41991;
squeal_samples[33187]=36840;
squeal_samples[33188]=32017;
squeal_samples[33189]=27507;
squeal_samples[33190]=23279;
squeal_samples[33191]=19336;
squeal_samples[33192]=15633;
squeal_samples[33193]=12178;
squeal_samples[33194]=8933;
squeal_samples[33195]=5905;
squeal_samples[33196]=4200;
squeal_samples[33197]=6770;
squeal_samples[33198]=9632;
squeal_samples[33199]=12368;
squeal_samples[33200]=14983;
squeal_samples[33201]=17482;
squeal_samples[33202]=19876;
squeal_samples[33203]=22156;
squeal_samples[33204]=24349;
squeal_samples[33205]=26427;
squeal_samples[33206]=28432;
squeal_samples[33207]=30326;
squeal_samples[33208]=32161;
squeal_samples[33209]=33887;
squeal_samples[33210]=35555;
squeal_samples[33211]=37139;
squeal_samples[33212]=38657;
squeal_samples[33213]=40103;
squeal_samples[33214]=41482;
squeal_samples[33215]=42807;
squeal_samples[33216]=44063;
squeal_samples[33217]=45270;
squeal_samples[33218]=46421;
squeal_samples[33219]=47514;
squeal_samples[33220]=48566;
squeal_samples[33221]=49562;
squeal_samples[33222]=50524;
squeal_samples[33223]=51438;
squeal_samples[33224]=52306;
squeal_samples[33225]=53146;
squeal_samples[33226]=53940;
squeal_samples[33227]=54490;
squeal_samples[33228]=50386;
squeal_samples[33229]=44703;
squeal_samples[33230]=39374;
squeal_samples[33231]=34395;
squeal_samples[33232]=29722;
squeal_samples[33233]=25361;
squeal_samples[33234]=21267;
squeal_samples[33235]=17455;
squeal_samples[33236]=13873;
squeal_samples[33237]=10522;
squeal_samples[33238]=7395;
squeal_samples[33239]=4503;
squeal_samples[33240]=5294;
squeal_samples[33241]=8206;
squeal_samples[33242]=11012;
squeal_samples[33243]=13684;
squeal_samples[33244]=16246;
squeal_samples[33245]=18686;
squeal_samples[33246]=21023;
squeal_samples[33247]=23258;
squeal_samples[33248]=25392;
squeal_samples[33249]=27432;
squeal_samples[33250]=29379;
squeal_samples[33251]=31248;
squeal_samples[33252]=33020;
squeal_samples[33253]=34727;
squeal_samples[33254]=36344;
squeal_samples[33255]=37903;
squeal_samples[33256]=39369;
squeal_samples[33257]=40796;
squeal_samples[33258]=42138;
squeal_samples[33259]=43435;
squeal_samples[33260]=44664;
squeal_samples[33261]=45836;
squeal_samples[33262]=46961;
squeal_samples[33263]=48036;
squeal_samples[33264]=49059;
squeal_samples[33265]=50041;
squeal_samples[33266]=50970;
squeal_samples[33267]=51867;
squeal_samples[33268]=52717;
squeal_samples[33269]=53536;
squeal_samples[33270]=54315;
squeal_samples[33271]=53151;
squeal_samples[33272]=47488;
squeal_samples[33273]=41985;
squeal_samples[33274]=36829;
squeal_samples[33275]=32009;
squeal_samples[33276]=27495;
squeal_samples[33277]=23270;
squeal_samples[33278]=19327;
squeal_samples[33279]=15615;
squeal_samples[33280]=12166;
squeal_samples[33281]=8913;
squeal_samples[33282]=5894;
squeal_samples[33283]=4176;
squeal_samples[33284]=6757;
squeal_samples[33285]=9615;
squeal_samples[33286]=12348;
squeal_samples[33287]=14966;
squeal_samples[33288]=17469;
squeal_samples[33289]=19852;
squeal_samples[33290]=22139;
squeal_samples[33291]=24324;
squeal_samples[33292]=26410;
squeal_samples[33293]=28407;
squeal_samples[33294]=30310;
squeal_samples[33295]=32135;
squeal_samples[33296]=33871;
squeal_samples[33297]=35530;
squeal_samples[33298]=37116;
squeal_samples[33299]=38634;
squeal_samples[33300]=40077;
squeal_samples[33301]=41462;
squeal_samples[33302]=42779;
squeal_samples[33303]=44044;
squeal_samples[33304]=45243;
squeal_samples[33305]=46393;
squeal_samples[33306]=47490;
squeal_samples[33307]=48542;
squeal_samples[33308]=49543;
squeal_samples[33309]=50498;
squeal_samples[33310]=51409;
squeal_samples[33311]=52289;
squeal_samples[33312]=53114;
squeal_samples[33313]=53919;
squeal_samples[33314]=54465;
squeal_samples[33315]=50367;
squeal_samples[33316]=44675;
squeal_samples[33317]=39355;
squeal_samples[33318]=34365;
squeal_samples[33319]=29705;
squeal_samples[33320]=25332;
squeal_samples[33321]=21247;
squeal_samples[33322]=17426;
squeal_samples[33323]=13848;
squeal_samples[33324]=10498;
squeal_samples[33325]=7371;
squeal_samples[33326]=4612;
squeal_samples[33327]=5970;
squeal_samples[33328]=8863;
squeal_samples[33329]=11632;
squeal_samples[33330]=14280;
squeal_samples[33331]=16810;
squeal_samples[33332]=19229;
squeal_samples[33333]=21540;
squeal_samples[33334]=23746;
squeal_samples[33335]=25860;
squeal_samples[33336]=27876;
squeal_samples[33337]=29811;
squeal_samples[33338]=31647;
squeal_samples[33339]=33414;
squeal_samples[33340]=35089;
squeal_samples[33341]=36694;
squeal_samples[33342]=38232;
squeal_samples[33343]=39693;
squeal_samples[33344]=41097;
squeal_samples[33345]=42429;
squeal_samples[33346]=43706;
squeal_samples[33347]=44919;
squeal_samples[33348]=46089;
squeal_samples[33349]=47191;
squeal_samples[33350]=48263;
squeal_samples[33351]=49269;
squeal_samples[33352]=50244;
squeal_samples[33353]=51161;
squeal_samples[33354]=52046;
squeal_samples[33355]=52893;
squeal_samples[33356]=53700;
squeal_samples[33357]=54468;
squeal_samples[33358]=51828;
squeal_samples[33359]=46041;
squeal_samples[33360]=40629;
squeal_samples[33361]=35559;
squeal_samples[33362]=30820;
squeal_samples[33363]=26376;
squeal_samples[33364]=22226;
squeal_samples[33365]=18338;
squeal_samples[33366]=14706;
squeal_samples[33367]=11295;
squeal_samples[33368]=8116;
squeal_samples[33369]=5128;
squeal_samples[33370]=5211;
squeal_samples[33371]=8139;
squeal_samples[33372]=10933;
squeal_samples[33373]=13617;
squeal_samples[33374]=16171;
squeal_samples[33375]=18620;
squeal_samples[33376]=20956;
squeal_samples[33377]=23191;
squeal_samples[33378]=25325;
squeal_samples[33379]=27370;
squeal_samples[33380]=29321;
squeal_samples[33381]=31177;
squeal_samples[33382]=32962;
squeal_samples[33383]=34663;
squeal_samples[33384]=36285;
squeal_samples[33385]=37839;
squeal_samples[33386]=39317;
squeal_samples[33387]=40736;
squeal_samples[33388]=42085;
squeal_samples[33389]=43378;
squeal_samples[33390]=44609;
squeal_samples[33391]=45784;
squeal_samples[33392]=46913;
squeal_samples[33393]=47982;
squeal_samples[33394]=49008;
squeal_samples[33395]=49986;
squeal_samples[33396]=50924;
squeal_samples[33397]=51813;
squeal_samples[33398]=52667;
squeal_samples[33399]=53487;
squeal_samples[33400]=54263;
squeal_samples[33401]=53103;
squeal_samples[33402]=47435;
squeal_samples[33403]=41936;
squeal_samples[33404]=36783;
squeal_samples[33405]=31965;
squeal_samples[33406]=27449;
squeal_samples[33407]=23227;
squeal_samples[33408]=19277;
squeal_samples[33409]=15577;
squeal_samples[33410]=12113;
squeal_samples[33411]=8880;
squeal_samples[33412]=5844;
squeal_samples[33413]=4627;
squeal_samples[33414]=7401;
squeal_samples[33415]=10234;
squeal_samples[33416]=12937;
squeal_samples[33417]=15530;
squeal_samples[33418]=18004;
squeal_samples[33419]=20368;
squeal_samples[33420]=22623;
squeal_samples[33421]=24788;
squeal_samples[33422]=26850;
squeal_samples[33423]=28830;
squeal_samples[33424]=30711;
squeal_samples[33425]=32512;
squeal_samples[33426]=34233;
squeal_samples[33427]=35877;
squeal_samples[33428]=37445;
squeal_samples[33429]=38942;
squeal_samples[33430]=40374;
squeal_samples[33431]=41743;
squeal_samples[33432]=43042;
squeal_samples[33433]=44294;
squeal_samples[33434]=45479;
squeal_samples[33435]=46621;
squeal_samples[33436]=47705;
squeal_samples[33437]=48743;
squeal_samples[33438]=49730;
squeal_samples[33439]=50681;
squeal_samples[33440]=51586;
squeal_samples[33441]=52444;
squeal_samples[33442]=53275;
squeal_samples[33443]=54057;
squeal_samples[33444]=53964;
squeal_samples[33445]=48859;
squeal_samples[33446]=43262;
squeal_samples[33447]=38027;
squeal_samples[33448]=33123;
squeal_samples[33449]=28534;
squeal_samples[33450]=24239;
squeal_samples[33451]=20222;
squeal_samples[33452]=16462;
squeal_samples[33453]=12945;
squeal_samples[33454]=9653;
squeal_samples[33455]=6570;
squeal_samples[33456]=4414;
squeal_samples[33457]=6664;
squeal_samples[33458]=9525;
squeal_samples[33459]=12263;
squeal_samples[33460]=14879;
squeal_samples[33461]=17386;
squeal_samples[33462]=19769;
squeal_samples[33463]=22063;
squeal_samples[33464]=24242;
squeal_samples[33465]=26332;
squeal_samples[33466]=28325;
squeal_samples[33467]=30238;
squeal_samples[33468]=32054;
squeal_samples[33469]=33798;
squeal_samples[33470]=35455;
squeal_samples[33471]=37047;
squeal_samples[33472]=38561;
squeal_samples[33473]=40008;
squeal_samples[33474]=41392;
squeal_samples[33475]=42713;
squeal_samples[33476]=43972;
squeal_samples[33477]=45183;
squeal_samples[33478]=46322;
squeal_samples[33479]=47428;
squeal_samples[33480]=48474;
squeal_samples[33481]=49478;
squeal_samples[33482]=50437;
squeal_samples[33483]=51343;
squeal_samples[33484]=52228;
squeal_samples[33485]=53050;
squeal_samples[33486]=53855;
squeal_samples[33487]=54559;
squeal_samples[33488]=51130;
squeal_samples[33489]=45390;
squeal_samples[33490]=40012;
squeal_samples[33491]=34983;
squeal_samples[33492]=30276;
squeal_samples[33493]=25871;
squeal_samples[33494]=21746;
squeal_samples[33495]=17888;
squeal_samples[33496]=14280;
squeal_samples[33497]=10893;
squeal_samples[33498]=7736;
squeal_samples[33499]=4773;
squeal_samples[33500]=4875;
squeal_samples[33501]=7811;
squeal_samples[33502]=10618;
squeal_samples[33503]=13312;
squeal_samples[33504]=15882;
squeal_samples[33505]=18338;
squeal_samples[33506]=20683;
squeal_samples[33507]=22929;
squeal_samples[33508]=25080;
squeal_samples[33509]=27130;
squeal_samples[33510]=29092;
squeal_samples[33511]=30959;
squeal_samples[33512]=32751;
squeal_samples[33513]=34453;
squeal_samples[33514]=36092;
squeal_samples[33515]=37645;
squeal_samples[33516]=39133;
squeal_samples[33517]=40556;
squeal_samples[33518]=41916;
squeal_samples[33519]=43208;
squeal_samples[33520]=44451;
squeal_samples[33521]=45631;
squeal_samples[33522]=46765;
squeal_samples[33523]=47835;
squeal_samples[33524]=48870;
squeal_samples[33525]=49850;
squeal_samples[33526]=50791;
squeal_samples[33527]=51688;
squeal_samples[33528]=52547;
squeal_samples[33529]=53364;
squeal_samples[33530]=54149;
squeal_samples[33531]=53568;
squeal_samples[33532]=48130;
squeal_samples[33533]=42581;
squeal_samples[33534]=37385;
squeal_samples[33535]=32523;
squeal_samples[33536]=27969;
squeal_samples[33537]=23710;
squeal_samples[33538]=19721;
squeal_samples[33539]=15998;
squeal_samples[33540]=12505;
squeal_samples[33541]=9241;
squeal_samples[33542]=6181;
squeal_samples[33543]=4452;
squeal_samples[33544]=7008;
squeal_samples[33545]=9858;
squeal_samples[33546]=12577;
squeal_samples[33547]=15182;
squeal_samples[33548]=17665;
squeal_samples[33549]=20042;
squeal_samples[33550]=22313;
squeal_samples[33551]=24492;
squeal_samples[33552]=26563;
squeal_samples[33553]=28551;
squeal_samples[33554]=30443;
squeal_samples[33555]=32258;
squeal_samples[33556]=33986;
squeal_samples[33557]=35638;
squeal_samples[33558]=37216;
squeal_samples[33559]=38723;
squeal_samples[33560]=40162;
squeal_samples[33561]=41540;
squeal_samples[33562]=42847;
squeal_samples[33563]=44108;
squeal_samples[33564]=45298;
squeal_samples[33565]=46447;
squeal_samples[33566]=47534;
squeal_samples[33567]=48580;
squeal_samples[33568]=49577;
squeal_samples[33569]=50528;
squeal_samples[33570]=51435;
squeal_samples[33571]=52305;
squeal_samples[33572]=53133;
squeal_samples[33573]=53928;
squeal_samples[33574]=54471;
squeal_samples[33575]=50369;
squeal_samples[33576]=44673;
squeal_samples[33577]=39346;
squeal_samples[33578]=34355;
squeal_samples[33579]=29682;
squeal_samples[33580]=25315;
squeal_samples[33581]=21224;
squeal_samples[33582]=17401;
squeal_samples[33583]=13819;
squeal_samples[33584]=10465;
squeal_samples[33585]=7325;
squeal_samples[33586]=4577;
squeal_samples[33587]=5927;
squeal_samples[33588]=8823;
squeal_samples[33589]=11589;
squeal_samples[33590]=14230;
squeal_samples[33591]=16767;
squeal_samples[33592]=19177;
squeal_samples[33593]=21489;
squeal_samples[33594]=23695;
squeal_samples[33595]=25809;
squeal_samples[33596]=27824;
squeal_samples[33597]=29756;
squeal_samples[33598]=31590;
squeal_samples[33599]=33352;
squeal_samples[33600]=35032;
squeal_samples[33601]=36638;
squeal_samples[33602]=38169;
squeal_samples[33603]=39634;
squeal_samples[33604]=41033;
squeal_samples[33605]=42366;
squeal_samples[33606]=43646;
squeal_samples[33607]=44855;
squeal_samples[33608]=46023;
squeal_samples[33609]=47131;
squeal_samples[33610]=48190;
squeal_samples[33611]=49208;
squeal_samples[33612]=50170;
squeal_samples[33613]=51099;
squeal_samples[33614]=51975;
squeal_samples[33615]=52821;
squeal_samples[33616]=53627;
squeal_samples[33617]=54400;
squeal_samples[33618]=52542;
squeal_samples[33619]=46757;
squeal_samples[33620]=41294;
squeal_samples[33621]=36183;
squeal_samples[33622]=31390;
squeal_samples[33623]=26916;
squeal_samples[33624]=22713;
squeal_samples[33625]=18797;
squeal_samples[33626]=15123;
squeal_samples[33627]=11687;
squeal_samples[33628]=8469;
squeal_samples[33629]=5468;
squeal_samples[33630]=4846;
squeal_samples[33631]=7747;
squeal_samples[33632]=10551;
squeal_samples[33633]=13244;
squeal_samples[33634]=15816;
squeal_samples[33635]=18278;
squeal_samples[33636]=20621;
squeal_samples[33637]=22869;
squeal_samples[33638]=25018;
squeal_samples[33639]=27071;
squeal_samples[33640]=29029;
squeal_samples[33641]=30901;
squeal_samples[33642]=32692;
squeal_samples[33643]=34401;
squeal_samples[33644]=36034;
squeal_samples[33645]=37592;
squeal_samples[33646]=39082;
squeal_samples[33647]=40506;
squeal_samples[33648]=41862;
squeal_samples[33649]=43156;
squeal_samples[33650]=44398;
squeal_samples[33651]=45575;
squeal_samples[33652]=46715;
squeal_samples[33653]=47786;
squeal_samples[33654]=48818;
squeal_samples[33655]=49804;
squeal_samples[33656]=50737;
squeal_samples[33657]=51647;
squeal_samples[33658]=52495;
squeal_samples[33659]=53319;
squeal_samples[33660]=54106;
squeal_samples[33661]=53999;
squeal_samples[33662]=48892;
squeal_samples[33663]=43290;
squeal_samples[33664]=38049;
squeal_samples[33665]=33138;
squeal_samples[33666]=28547;
squeal_samples[33667]=24243;
squeal_samples[33668]=20223;
squeal_samples[33669]=16457;
squeal_samples[33670]=12940;
squeal_samples[33671]=9641;
squeal_samples[33672]=6556;
squeal_samples[33673]=4391;
squeal_samples[33674]=6643;
squeal_samples[33675]=9504;
squeal_samples[33676]=12234;
squeal_samples[33677]=14855;
squeal_samples[33678]=17357;
squeal_samples[33679]=19739;
squeal_samples[33680]=22028;
squeal_samples[33681]=24211;
squeal_samples[33682]=26298;
squeal_samples[33683]=28296;
squeal_samples[33684]=30197;
squeal_samples[33685]=32019;
squeal_samples[33686]=33758;
squeal_samples[33687]=35419;
squeal_samples[33688]=37003;
squeal_samples[33689]=38518;
squeal_samples[33690]=39964;
squeal_samples[33691]=41352;
squeal_samples[33692]=42665;
squeal_samples[33693]=43928;
squeal_samples[33694]=45131;
squeal_samples[33695]=46281;
squeal_samples[33696]=47379;
squeal_samples[33697]=48425;
squeal_samples[33698]=49425;
squeal_samples[33699]=50381;
squeal_samples[33700]=51298;
squeal_samples[33701]=52170;
squeal_samples[33702]=53000;
squeal_samples[33703]=53804;
squeal_samples[33704]=54507;
squeal_samples[33705]=51075;
squeal_samples[33706]=45330;
squeal_samples[33707]=39959;
squeal_samples[33708]=34929;
squeal_samples[33709]=30222;
squeal_samples[33710]=25812;
squeal_samples[33711]=21685;
squeal_samples[33712]=17830;
squeal_samples[33713]=14220;
squeal_samples[33714]=10832;
squeal_samples[33715]=7678;
squeal_samples[33716]=4754;
squeal_samples[33717]=5530;
squeal_samples[33718]=8429;
squeal_samples[33719]=11212;
squeal_samples[33720]=13875;
squeal_samples[33721]=16415;
squeal_samples[33722]=18848;
squeal_samples[33723]=21167;
squeal_samples[33724]=23392;
squeal_samples[33725]=25513;
squeal_samples[33726]=27544;
squeal_samples[33727]=29481;
squeal_samples[33728]=31332;
squeal_samples[33729]=33100;
squeal_samples[33730]=34794;
squeal_samples[33731]=36403;
squeal_samples[33732]=37947;
squeal_samples[33733]=39415;
squeal_samples[33734]=40822;
squeal_samples[33735]=42166;
squeal_samples[33736]=43448;
squeal_samples[33737]=44672;
squeal_samples[33738]=45841;
squeal_samples[33739]=46959;
squeal_samples[33740]=48026;
squeal_samples[33741]=49045;
squeal_samples[33742]=50012;
squeal_samples[33743]=50945;
squeal_samples[33744]=51836;
squeal_samples[33745]=52682;
squeal_samples[33746]=53497;
squeal_samples[33747]=54269;
squeal_samples[33748]=53101;
squeal_samples[33749]=47430;
squeal_samples[33750]=41925;
squeal_samples[33751]=36760;
squeal_samples[33752]=31940;
squeal_samples[33753]=27412;
squeal_samples[33754]=23192;
squeal_samples[33755]=19232;
squeal_samples[33756]=15533;
squeal_samples[33757]=12065;
squeal_samples[33758]=8824;
squeal_samples[33759]=5789;
squeal_samples[33760]=4575;
squeal_samples[33761]=7339;
squeal_samples[33762]=10174;
squeal_samples[33763]=12878;
squeal_samples[33764]=15463;
squeal_samples[33765]=17941;
squeal_samples[33766]=20295;
squeal_samples[33767]=22554;
squeal_samples[33768]=24715;
squeal_samples[33769]=26781;
squeal_samples[33770]=28753;
squeal_samples[33771]=30635;
squeal_samples[33772]=32436;
squeal_samples[33773]=34152;
squeal_samples[33774]=35795;
squeal_samples[33775]=37362;
squeal_samples[33776]=38862;
squeal_samples[33777]=40293;
squeal_samples[33778]=41654;
squeal_samples[33779]=42963;
squeal_samples[33780]=44205;
squeal_samples[33781]=45398;
squeal_samples[33782]=46535;
squeal_samples[33783]=47616;
squeal_samples[33784]=48657;
squeal_samples[33785]=49643;
squeal_samples[33786]=50590;
squeal_samples[33787]=51490;
squeal_samples[33788]=52355;
squeal_samples[33789]=53184;
squeal_samples[33790]=53966;
squeal_samples[33791]=54247;
squeal_samples[33792]=49575;
squeal_samples[33793]=43931;
squeal_samples[33794]=38646;
squeal_samples[33795]=33698;
squeal_samples[33796]=29066;
squeal_samples[33797]=24730;
squeal_samples[33798]=20670;
squeal_samples[33799]=16882;
squeal_samples[33800]=13325;
squeal_samples[33801]=9999;
squeal_samples[33802]=6895;
squeal_samples[33803]=4388;
squeal_samples[33804]=6239;
squeal_samples[33805]=9107;
squeal_samples[33806]=11870;
squeal_samples[33807]=14493;
squeal_samples[33808]=17010;
squeal_samples[33809]=19410;
squeal_samples[33810]=21710;
squeal_samples[33811]=23904;
squeal_samples[33812]=26004;
squeal_samples[33813]=28012;
squeal_samples[33814]=29929;
squeal_samples[33815]=31756;
squeal_samples[33816]=33503;
squeal_samples[33817]=35177;
squeal_samples[33818]=36766;
squeal_samples[33819]=38299;
squeal_samples[33820]=39745;
squeal_samples[33821]=41140;
squeal_samples[33822]=42466;
squeal_samples[33823]=43736;
squeal_samples[33824]=44947;
squeal_samples[33825]=46103;
squeal_samples[33826]=47203;
squeal_samples[33827]=48259;
squeal_samples[33828]=49265;
squeal_samples[33829]=50230;
squeal_samples[33830]=51145;
squeal_samples[33831]=52023;
squeal_samples[33832]=52864;
squeal_samples[33833]=53666;
squeal_samples[33834]=54431;
squeal_samples[33835]=52568;
squeal_samples[33836]=46777;
squeal_samples[33837]=41310;
squeal_samples[33838]=36190;
squeal_samples[33839]=31400;
squeal_samples[33840]=26915;
squeal_samples[33841]=22711;
squeal_samples[33842]=18791;
squeal_samples[33843]=15117;
squeal_samples[33844]=11670;
squeal_samples[33845]=8459;
squeal_samples[33846]=5443;
squeal_samples[33847]=4244;
squeal_samples[33848]=7029;
squeal_samples[33849]=9870;
squeal_samples[33850]=12588;
squeal_samples[33851]=15183;
squeal_samples[33852]=17671;
squeal_samples[33853]=20037;
squeal_samples[33854]=22312;
squeal_samples[33855]=24477;
squeal_samples[33856]=26552;
squeal_samples[33857]=28530;
squeal_samples[33858]=30428;
squeal_samples[33859]=32229;
squeal_samples[33860]=33960;
squeal_samples[33861]=35607;
squeal_samples[33862]=37185;
squeal_samples[33863]=38691;
squeal_samples[33864]=40124;
squeal_samples[33865]=41502;
squeal_samples[33866]=42806;
squeal_samples[33867]=44059;
squeal_samples[33868]=45257;
squeal_samples[33869]=46396;
squeal_samples[33870]=47487;
squeal_samples[33871]=48527;
squeal_samples[33872]=49520;
squeal_samples[33873]=50472;
squeal_samples[33874]=51377;
squeal_samples[33875]=52245;
squeal_samples[33876]=53073;
squeal_samples[33877]=53869;
squeal_samples[33878]=54568;
squeal_samples[33879]=51129;
squeal_samples[33880]=45379;
squeal_samples[33881]=39998;
squeal_samples[33882]=34967;
squeal_samples[33883]=30246;
squeal_samples[33884]=25837;
squeal_samples[33885]=21708;
squeal_samples[33886]=17842;
squeal_samples[33887]=14231;
squeal_samples[33888]=10842;
squeal_samples[33889]=7680;
squeal_samples[33890]=4713;
squeal_samples[33891]=4808;
squeal_samples[33892]=7744;
squeal_samples[33893]=10554;
squeal_samples[33894]=13243;
squeal_samples[33895]=15812;
squeal_samples[33896]=18265;
squeal_samples[33897]=20611;
squeal_samples[33898]=22853;
squeal_samples[33899]=24997;
squeal_samples[33900]=27048;
squeal_samples[33901]=29008;
squeal_samples[33902]=30879;
squeal_samples[33903]=32665;
squeal_samples[33904]=34367;
squeal_samples[33905]=36003;
squeal_samples[33906]=37557;
squeal_samples[33907]=39048;
squeal_samples[33908]=40464;
squeal_samples[33909]=41825;
squeal_samples[33910]=43118;
squeal_samples[33911]=44358;
squeal_samples[33912]=45534;
squeal_samples[33913]=46664;
squeal_samples[33914]=47744;
squeal_samples[33915]=48768;
squeal_samples[33916]=49754;
squeal_samples[33917]=50690;
squeal_samples[33918]=51590;
squeal_samples[33919]=52448;
squeal_samples[33920]=53264;
squeal_samples[33921]=54050;
squeal_samples[33922]=54314;
squeal_samples[33923]=49648;
squeal_samples[33924]=43990;
squeal_samples[33925]=38701;
squeal_samples[33926]=33741;
squeal_samples[33927]=29106;
squeal_samples[33928]=24764;
squeal_samples[33929]=20706;
squeal_samples[33930]=16909;
squeal_samples[33931]=13350;
squeal_samples[33932]=10025;
squeal_samples[33933]=6906;
squeal_samples[33934]=4404;
squeal_samples[33935]=6246;
squeal_samples[33936]=9121;
squeal_samples[33937]=11874;
squeal_samples[33938]=14499;
squeal_samples[33939]=17016;
squeal_samples[33940]=19409;
squeal_samples[33941]=21705;
squeal_samples[33942]=23905;
squeal_samples[33943]=25999;
squeal_samples[33944]=28006;
squeal_samples[33945]=29919;
squeal_samples[33946]=31749;
squeal_samples[33947]=33500;
squeal_samples[33948]=35164;
squeal_samples[33949]=36758;
squeal_samples[33950]=38287;
squeal_samples[33951]=39735;
squeal_samples[33952]=41123;
squeal_samples[33953]=42450;
squeal_samples[33954]=43716;
squeal_samples[33955]=44925;
squeal_samples[33956]=46081;
squeal_samples[33957]=47182;
squeal_samples[33958]=48237;
squeal_samples[33959]=49245;
squeal_samples[33960]=50208;
squeal_samples[33961]=51124;
squeal_samples[33962]=52000;
squeal_samples[33963]=52839;
squeal_samples[33964]=53638;
squeal_samples[33965]=54405;
squeal_samples[33966]=52541;
squeal_samples[33967]=46749;
squeal_samples[33968]=41284;
squeal_samples[33969]=36163;
squeal_samples[33970]=31367;
squeal_samples[33971]=26882;
squeal_samples[33972]=22685;
squeal_samples[33973]=18759;
squeal_samples[33974]=15083;
squeal_samples[33975]=11639;
squeal_samples[33976]=8423;
squeal_samples[33977]=5413;
squeal_samples[33978]=4791;
squeal_samples[33979]=7687;
squeal_samples[33980]=10496;
squeal_samples[33981]=13183;
squeal_samples[33982]=15756;
squeal_samples[33983]=18212;
squeal_samples[33984]=20558;
squeal_samples[33985]=22803;
squeal_samples[33986]=24948;
squeal_samples[33987]=27003;
squeal_samples[33988]=28960;
squeal_samples[33989]=30833;
squeal_samples[33990]=32617;
squeal_samples[33991]=34329;
squeal_samples[33992]=35953;
squeal_samples[33993]=37519;
squeal_samples[33994]=39003;
squeal_samples[33995]=40426;
squeal_samples[33996]=41782;
squeal_samples[33997]=43079;
squeal_samples[33998]=44315;
squeal_samples[33999]=45500;
squeal_samples[34000]=46627;
squeal_samples[34001]=47703;
squeal_samples[34002]=48734;
squeal_samples[34003]=49715;
squeal_samples[34004]=50659;
squeal_samples[34005]=51550;
squeal_samples[34006]=52415;
squeal_samples[34007]=53227;
squeal_samples[34008]=54014;
squeal_samples[34009]=54280;
squeal_samples[34010]=49610;
squeal_samples[34011]=43962;
squeal_samples[34012]=38664;
squeal_samples[34013]=33712;
squeal_samples[34014]=29073;
squeal_samples[34015]=24738;
squeal_samples[34016]=20672;
squeal_samples[34017]=16881;
squeal_samples[34018]=13321;
squeal_samples[34019]=9991;
squeal_samples[34020]=6881;
squeal_samples[34021]=4369;
squeal_samples[34022]=6223;
squeal_samples[34023]=9093;
squeal_samples[34024]=11841;
squeal_samples[34025]=14471;
squeal_samples[34026]=16984;
squeal_samples[34027]=19386;
squeal_samples[34028]=21679;
squeal_samples[34029]=23877;
squeal_samples[34030]=25971;
squeal_samples[34031]=27980;
squeal_samples[34032]=29891;
squeal_samples[34033]=31722;
squeal_samples[34034]=33467;
squeal_samples[34035]=35142;
squeal_samples[34036]=36732;
squeal_samples[34037]=38257;
squeal_samples[34038]=39706;
squeal_samples[34039]=41097;
squeal_samples[34040]=42428;
squeal_samples[34041]=43688;
squeal_samples[34042]=44902;
squeal_samples[34043]=46056;
squeal_samples[34044]=47158;
squeal_samples[34045]=48212;
squeal_samples[34046]=49221;
squeal_samples[34047]=50176;
squeal_samples[34048]=51096;
squeal_samples[34049]=51976;
squeal_samples[34050]=52812;
squeal_samples[34051]=53616;
squeal_samples[34052]=54377;
squeal_samples[34053]=52520;
squeal_samples[34054]=46723;
squeal_samples[34055]=41254;
squeal_samples[34056]=36139;
squeal_samples[34057]=31342;
squeal_samples[34058]=26858;
squeal_samples[34059]=22661;
squeal_samples[34060]=18732;
squeal_samples[34061]=15061;
squeal_samples[34062]=11613;
squeal_samples[34063]=8401;
squeal_samples[34064]=5381;
squeal_samples[34065]=4768;
squeal_samples[34066]=7662;
squeal_samples[34067]=10469;
squeal_samples[34068]=13165;
squeal_samples[34069]=15724;
squeal_samples[34070]=18193;
squeal_samples[34071]=20532;
squeal_samples[34072]=22777;
squeal_samples[34073]=24926;
squeal_samples[34074]=26977;
squeal_samples[34075]=28935;
squeal_samples[34076]=30804;
squeal_samples[34077]=32592;
squeal_samples[34078]=34305;
squeal_samples[34079]=35929;
squeal_samples[34080]=37489;
squeal_samples[34081]=38977;
squeal_samples[34082]=40404;
squeal_samples[34083]=41754;
squeal_samples[34084]=43059;
squeal_samples[34085]=44288;
squeal_samples[34086]=45476;
squeal_samples[34087]=46603;
squeal_samples[34088]=47678;
squeal_samples[34089]=48709;
squeal_samples[34090]=49693;
squeal_samples[34091]=50632;
squeal_samples[34092]=51527;
squeal_samples[34093]=52391;
squeal_samples[34094]=53201;
squeal_samples[34095]=53991;
squeal_samples[34096]=54256;
squeal_samples[34097]=49584;
squeal_samples[34098]=43940;
squeal_samples[34099]=38637;
squeal_samples[34100]=33689;
squeal_samples[34101]=29050;
squeal_samples[34102]=24711;
squeal_samples[34103]=20651;
squeal_samples[34104]=16853;
squeal_samples[34105]=13299;
squeal_samples[34106]=9966;
squeal_samples[34107]=6856;
squeal_samples[34108]=4347;
squeal_samples[34109]=6196;
squeal_samples[34110]=9071;
squeal_samples[34111]=11815;
squeal_samples[34112]=14448;
squeal_samples[34113]=16959;
squeal_samples[34114]=19362;
squeal_samples[34115]=21656;
squeal_samples[34116]=23850;
squeal_samples[34117]=25950;
squeal_samples[34118]=27952;
squeal_samples[34119]=29870;
squeal_samples[34120]=31696;
squeal_samples[34121]=33444;
squeal_samples[34122]=35116;
squeal_samples[34123]=36710;
squeal_samples[34124]=38231;
squeal_samples[34125]=39682;
squeal_samples[34126]=41074;
squeal_samples[34127]=42402;
squeal_samples[34128]=43665;
squeal_samples[34129]=44879;
squeal_samples[34130]=46029;
squeal_samples[34131]=47137;
squeal_samples[34132]=48185;
squeal_samples[34133]=49198;
squeal_samples[34134]=50152;
squeal_samples[34135]=51071;
squeal_samples[34136]=51952;
squeal_samples[34137]=52789;
squeal_samples[34138]=53590;
squeal_samples[34139]=54356;
squeal_samples[34140]=52491;
squeal_samples[34141]=46703;
squeal_samples[34142]=41228;
squeal_samples[34143]=36115;
squeal_samples[34144]=31319;
squeal_samples[34145]=26832;
squeal_samples[34146]=22637;
squeal_samples[34147]=18710;
squeal_samples[34148]=15035;
squeal_samples[34149]=11590;
squeal_samples[34150]=8375;
squeal_samples[34151]=5358;
squeal_samples[34152]=4744;
squeal_samples[34153]=7637;
squeal_samples[34154]=10448;
squeal_samples[34155]=13135;
squeal_samples[34156]=15706;
squeal_samples[34157]=18164;
squeal_samples[34158]=20511;
squeal_samples[34159]=22752;
squeal_samples[34160]=24901;
squeal_samples[34161]=26953;
squeal_samples[34162]=28912;
squeal_samples[34163]=30779;
squeal_samples[34164]=32570;
squeal_samples[34165]=34277;
squeal_samples[34166]=35909;
squeal_samples[34167]=37460;
squeal_samples[34168]=38959;
squeal_samples[34169]=40374;
squeal_samples[34170]=41735;
squeal_samples[34171]=43030;
squeal_samples[34172]=44267;
squeal_samples[34173]=45451;
squeal_samples[34174]=46578;
squeal_samples[34175]=47655;
squeal_samples[34176]=48683;
squeal_samples[34177]=49671;
squeal_samples[34178]=50606;
squeal_samples[34179]=51505;
squeal_samples[34180]=52364;
squeal_samples[34181]=53177;
squeal_samples[34182]=53969;
squeal_samples[34183]=54499;
squeal_samples[34184]=50385;
squeal_samples[34185]=44678;
squeal_samples[34186]=39331;
squeal_samples[34187]=34340;
squeal_samples[34188]=29653;
squeal_samples[34189]=25276;
squeal_samples[34190]=21173;
squeal_samples[34191]=17346;
squeal_samples[34192]=13757;
squeal_samples[34193]=10395;
squeal_samples[34194]=7254;
squeal_samples[34195]=4492;
squeal_samples[34196]=5841;
squeal_samples[34197]=8730;
squeal_samples[34198]=11493;
squeal_samples[34199]=14137;
squeal_samples[34200]=16656;
squeal_samples[34201]=19079;
squeal_samples[34202]=21377;
squeal_samples[34203]=23585;
squeal_samples[34204]=25696;
squeal_samples[34205]=27707;
squeal_samples[34206]=29638;
squeal_samples[34207]=31468;
squeal_samples[34208]=33233;
squeal_samples[34209]=34905;
squeal_samples[34210]=36508;
squeal_samples[34211]=38038;
squeal_samples[34212]=39502;
squeal_samples[34213]=40897;
squeal_samples[34214]=42232;
squeal_samples[34215]=43505;
squeal_samples[34216]=44724;
squeal_samples[34217]=45882;
squeal_samples[34218]=46991;
squeal_samples[34219]=48049;
squeal_samples[34220]=49058;
squeal_samples[34221]=50027;
squeal_samples[34222]=50947;
squeal_samples[34223]=51831;
squeal_samples[34224]=52671;
squeal_samples[34225]=53479;
squeal_samples[34226]=54248;
squeal_samples[34227]=53654;
squeal_samples[34228]=48197;
squeal_samples[34229]=42631;
squeal_samples[34230]=37417;
squeal_samples[34231]=32542;
squeal_samples[34232]=27973;
squeal_samples[34233]=23707;
squeal_samples[34234]=19699;
squeal_samples[34235]=15969;
squeal_samples[34236]=12460;
squeal_samples[34237]=9189;
squeal_samples[34238]=6117;
squeal_samples[34239]=4375;
squeal_samples[34240]=6938;
squeal_samples[34241]=9767;
squeal_samples[34242]=12490;
squeal_samples[34243]=15088;
squeal_samples[34244]=17572;
squeal_samples[34245]=19943;
squeal_samples[34246]=22213;
squeal_samples[34247]=24377;
squeal_samples[34248]=26454;
squeal_samples[34249]=28430;
squeal_samples[34250]=30328;
squeal_samples[34251]=32131;
squeal_samples[34252]=33862;
squeal_samples[34253]=35504;
squeal_samples[34254]=37086;
squeal_samples[34255]=38580;
squeal_samples[34256]=40026;
squeal_samples[34257]=41393;
squeal_samples[34258]=42703;
squeal_samples[34259]=43956;
squeal_samples[34260]=45150;
squeal_samples[34261]=46295;
squeal_samples[34262]=47380;
squeal_samples[34263]=48424;
squeal_samples[34264]=49414;
squeal_samples[34265]=50369;
squeal_samples[34266]=51273;
squeal_samples[34267]=52138;
squeal_samples[34268]=52967;
squeal_samples[34269]=53760;
squeal_samples[34270]=54514;
squeal_samples[34271]=51857;
squeal_samples[34272]=46054;
squeal_samples[34273]=40625;
squeal_samples[34274]=35539;
squeal_samples[34275]=30785;
squeal_samples[34276]=26322;
squeal_samples[34277]=22166;
squeal_samples[34278]=18256;
squeal_samples[34279]=14618;
squeal_samples[34280]=11193;
squeal_samples[34281]=8004;
squeal_samples[34282]=5006;
squeal_samples[34283]=5084;
squeal_samples[34284]=7997;
squeal_samples[34285]=10794;
squeal_samples[34286]=13463;
squeal_samples[34287]=16023;
squeal_samples[34288]=18466;
squeal_samples[34289]=20794;
squeal_samples[34290]=23026;
squeal_samples[34291]=25160;
squeal_samples[34292]=27193;
squeal_samples[34293]=29143;
squeal_samples[34294]=30998;
squeal_samples[34295]=32778;
squeal_samples[34296]=34476;
squeal_samples[34297]=36095;
squeal_samples[34298]=37642;
squeal_samples[34299]=39125;
squeal_samples[34300]=40527;
squeal_samples[34301]=41886;
squeal_samples[34302]=43166;
squeal_samples[34303]=44401;
squeal_samples[34304]=45573;
squeal_samples[34305]=46694;
squeal_samples[34306]=47767;
squeal_samples[34307]=48789;
squeal_samples[34308]=49770;
squeal_samples[34309]=50696;
squeal_samples[34310]=51595;
squeal_samples[34311]=52441;
squeal_samples[34312]=53259;
squeal_samples[34313]=54035;
squeal_samples[34314]=54296;
squeal_samples[34315]=49628;
squeal_samples[34316]=43962;
squeal_samples[34317]=38666;
squeal_samples[34318]=33713;
squeal_samples[34319]=29063;
squeal_samples[34320]=24726;
squeal_samples[34321]=20654;
squeal_samples[34322]=16855;
squeal_samples[34323]=13292;
squeal_samples[34324]=9963;
squeal_samples[34325]=6844;
squeal_samples[34326]=4336;
squeal_samples[34327]=6184;
squeal_samples[34328]=9049;
squeal_samples[34329]=11799;
squeal_samples[34330]=14423;
squeal_samples[34331]=16941;
squeal_samples[34332]=19332;
squeal_samples[34333]=21632;
squeal_samples[34334]=23821;
squeal_samples[34335]=25920;
squeal_samples[34336]=27920;
squeal_samples[34337]=29835;
squeal_samples[34338]=31667;
squeal_samples[34339]=33410;
squeal_samples[34340]=35080;
squeal_samples[34341]=36672;
squeal_samples[34342]=38192;
squeal_samples[34343]=39647;
squeal_samples[34344]=41035;
squeal_samples[34345]=42359;
squeal_samples[34346]=43624;
squeal_samples[34347]=44833;
squeal_samples[34348]=45989;
squeal_samples[34349]=47092;
squeal_samples[34350]=48143;
squeal_samples[34351]=49150;
squeal_samples[34352]=50109;
squeal_samples[34353]=51028;
squeal_samples[34354]=51903;
squeal_samples[34355]=52741;
squeal_samples[34356]=53541;
squeal_samples[34357]=54307;
squeal_samples[34358]=53123;
squeal_samples[34359]=47447;
squeal_samples[34360]=41925;
squeal_samples[34361]=36756;
squeal_samples[34362]=31916;
squeal_samples[34363]=27388;
squeal_samples[34364]=23153;
squeal_samples[34365]=19189;
squeal_samples[34366]=15480;
squeal_samples[34367]=12004;
squeal_samples[34368]=8757;
squeal_samples[34369]=5717;
squeal_samples[34370]=4495;
squeal_samples[34371]=7256;
squeal_samples[34372]=10087;
squeal_samples[34373]=12780;
squeal_samples[34374]=15375;
squeal_samples[34375]=17834;
squeal_samples[34376]=20201;
squeal_samples[34377]=22452;
squeal_samples[34378]=24611;
squeal_samples[34379]=26671;
squeal_samples[34380]=28641;
squeal_samples[34381]=30521;
squeal_samples[34382]=32313;
squeal_samples[34383]=34039;
squeal_samples[34384]=35671;
squeal_samples[34385]=37244;
squeal_samples[34386]=38733;
squeal_samples[34387]=40161;
squeal_samples[34388]=41529;
squeal_samples[34389]=42830;
squeal_samples[34390]=44074;
squeal_samples[34391]=45260;
squeal_samples[34392]=46398;
squeal_samples[34393]=47479;
squeal_samples[34394]=48515;
squeal_samples[34395]=49498;
squeal_samples[34396]=50449;
squeal_samples[34397]=51346;
squeal_samples[34398]=52214;
squeal_samples[34399]=53033;
squeal_samples[34400]=53820;
squeal_samples[34401]=54519;
squeal_samples[34402]=51074;
squeal_samples[34403]=45322;
squeal_samples[34404]=39935;
squeal_samples[34405]=34895;
squeal_samples[34406]=30171;
squeal_samples[34407]=25759;
squeal_samples[34408]=21621;
squeal_samples[34409]=17760;
squeal_samples[34410]=14138;
squeal_samples[34411]=10750;
squeal_samples[34412]=7581;
squeal_samples[34413]=4663;
squeal_samples[34414]=5418;
squeal_samples[34415]=8323;
squeal_samples[34416]=11099;
squeal_samples[34417]=13756;
squeal_samples[34418]=16298;
squeal_samples[34419]=18724;
squeal_samples[34420]=21042;
squeal_samples[34421]=23264;
squeal_samples[34422]=25377;
squeal_samples[34423]=27413;
squeal_samples[34424]=29337;
squeal_samples[34425]=31196;
squeal_samples[34426]=32957;
squeal_samples[34427]=34650;
squeal_samples[34428]=36259;
squeal_samples[34429]=37794;
squeal_samples[34430]=39266;
squeal_samples[34431]=40672;
squeal_samples[34432]=42008;
squeal_samples[34433]=43295;
squeal_samples[34434]=44507;
squeal_samples[34435]=45689;
squeal_samples[34436]=46793;
squeal_samples[34437]=47864;
squeal_samples[34438]=48878;
squeal_samples[34439]=49857;
squeal_samples[34440]=50774;
squeal_samples[34441]=51670;
squeal_samples[34442]=52510;
squeal_samples[34443]=53322;
squeal_samples[34444]=54098;
squeal_samples[34445]=53982;
squeal_samples[34446]=48862;
squeal_samples[34447]=43250;
squeal_samples[34448]=37993;
squeal_samples[34449]=33077;
squeal_samples[34450]=28474;
squeal_samples[34451]=24160;
squeal_samples[34452]=20134;
squeal_samples[34453]=16358;
squeal_samples[34454]=12829;
squeal_samples[34455]=9528;
squeal_samples[34456]=6431;
squeal_samples[34457]=4269;
squeal_samples[34458]=6507;
squeal_samples[34459]=9370;
squeal_samples[34460]=12096;
squeal_samples[34461]=14712;
squeal_samples[34462]=17209;
squeal_samples[34463]=19592;
squeal_samples[34464]=21873;
squeal_samples[34465]=24055;
squeal_samples[34466]=26138;
squeal_samples[34467]=28131;
squeal_samples[34468]=30035;
squeal_samples[34469]=31853;
squeal_samples[34470]=33590;
squeal_samples[34471]=35249;
squeal_samples[34472]=36834;
squeal_samples[34473]=38343;
squeal_samples[34474]=39791;
squeal_samples[34475]=41169;
squeal_samples[34476]=42488;
squeal_samples[34477]=43746;
squeal_samples[34478]=44946;
squeal_samples[34479]=46097;
squeal_samples[34480]=47191;
squeal_samples[34481]=48242;
squeal_samples[34482]=49238;
squeal_samples[34483]=50196;
squeal_samples[34484]=51102;
squeal_samples[34485]=51978;
squeal_samples[34486]=52810;
squeal_samples[34487]=53605;
squeal_samples[34488]=54365;
squeal_samples[34489]=52498;
squeal_samples[34490]=46699;
squeal_samples[34491]=41225;
squeal_samples[34492]=36100;
squeal_samples[34493]=31304;
squeal_samples[34494]=26808;
squeal_samples[34495]=22611;
squeal_samples[34496]=18674;
squeal_samples[34497]=15004;
squeal_samples[34498]=11549;
squeal_samples[34499]=8334;
squeal_samples[34500]=5310;
squeal_samples[34501]=4697;
squeal_samples[34502]=7586;
squeal_samples[34503]=10393;
squeal_samples[34504]=13082;
squeal_samples[34505]=15649;
squeal_samples[34506]=18105;
squeal_samples[34507]=20450;
squeal_samples[34508]=22691;
squeal_samples[34509]=24836;
squeal_samples[34510]=26888;
squeal_samples[34511]=28846;
squeal_samples[34512]=30713;
squeal_samples[34513]=32504;
squeal_samples[34514]=34206;
squeal_samples[34515]=35843;
squeal_samples[34516]=37397;
squeal_samples[34517]=38883;
squeal_samples[34518]=40303;
squeal_samples[34519]=41655;
squeal_samples[34520]=42955;
squeal_samples[34521]=44191;
squeal_samples[34522]=45372;
squeal_samples[34523]=46505;
squeal_samples[34524]=47575;
squeal_samples[34525]=48611;
squeal_samples[34526]=49591;
squeal_samples[34527]=50525;
squeal_samples[34528]=51425;
squeal_samples[34529]=52277;
squeal_samples[34530]=53102;
squeal_samples[34531]=53880;
squeal_samples[34532]=54578;
squeal_samples[34533]=51129;
squeal_samples[34534]=45366;
squeal_samples[34535]=39975;
squeal_samples[34536]=34927;
squeal_samples[34537]=30206;
squeal_samples[34538]=25782;
squeal_samples[34539]=21649;
squeal_samples[34540]=17778;
squeal_samples[34541]=14154;
squeal_samples[34542]=10765;
squeal_samples[34543]=7589;
squeal_samples[34544]=4669;
squeal_samples[34545]=5420;
squeal_samples[34546]=8329;
squeal_samples[34547]=11101;
squeal_samples[34548]=13762;
squeal_samples[34549]=16294;
squeal_samples[34550]=18725;
squeal_samples[34551]=21040;
squeal_samples[34552]=23256;
squeal_samples[34553]=25378;
squeal_samples[34554]=27403;
squeal_samples[34555]=29334;
squeal_samples[34556]=31185;
squeal_samples[34557]=32948;
squeal_samples[34558]=34636;
squeal_samples[34559]=36247;
squeal_samples[34560]=37783;
squeal_samples[34561]=39253;
squeal_samples[34562]=40653;
squeal_samples[34563]=41993;
squeal_samples[34564]=43273;
squeal_samples[34565]=44495;
squeal_samples[34566]=45661;
squeal_samples[34567]=46779;
squeal_samples[34568]=47843;
squeal_samples[34569]=48859;
squeal_samples[34570]=49829;
squeal_samples[34571]=50760;
squeal_samples[34572]=51644;
squeal_samples[34573]=52488;
squeal_samples[34574]=53300;
squeal_samples[34575]=54072;
squeal_samples[34576]=54329;
squeal_samples[34577]=49648;
squeal_samples[34578]=43983;
squeal_samples[34579]=38681;
squeal_samples[34580]=33716;
squeal_samples[34581]=29070;
squeal_samples[34582]=24718;
squeal_samples[34583]=20650;
squeal_samples[34584]=16843;
squeal_samples[34585]=13281;
squeal_samples[34586]=9942;
squeal_samples[34587]=6824;
squeal_samples[34588]=4315;
squeal_samples[34589]=6152;
squeal_samples[34590]=9028;
squeal_samples[34591]=11765;
squeal_samples[34592]=14401;
squeal_samples[34593]=16899;
squeal_samples[34594]=19300;
squeal_samples[34595]=21595;
squeal_samples[34596]=23786;
squeal_samples[34597]=25884;
squeal_samples[34598]=27884;
squeal_samples[34599]=29796;
squeal_samples[34600]=31623;
squeal_samples[34601]=33367;
squeal_samples[34602]=35036;
squeal_samples[34603]=36628;
squeal_samples[34604]=38145;
squeal_samples[34605]=39601;
squeal_samples[34606]=40987;
squeal_samples[34607]=42314;
squeal_samples[34608]=43577;
squeal_samples[34609]=44783;
squeal_samples[34610]=45936;
squeal_samples[34611]=47041;
squeal_samples[34612]=48090;
squeal_samples[34613]=49099;
squeal_samples[34614]=50057;
squeal_samples[34615]=50972;
squeal_samples[34616]=51845;
squeal_samples[34617]=52683;
squeal_samples[34618]=53485;
squeal_samples[34619]=54247;
squeal_samples[34620]=53651;
squeal_samples[34621]=48185;
squeal_samples[34622]=42614;
squeal_samples[34623]=37399;
squeal_samples[34624]=32516;
squeal_samples[34625]=27946;
squeal_samples[34626]=23664;
squeal_samples[34627]=19667;
squeal_samples[34628]=15920;
squeal_samples[34629]=12418;
squeal_samples[34630]=9130;
squeal_samples[34631]=6066;
squeal_samples[34632]=4321;
squeal_samples[34633]=6877;
squeal_samples[34634]=9710;
squeal_samples[34635]=12430;
squeal_samples[34636]=15024;
squeal_samples[34637]=17507;
squeal_samples[34638]=19872;
squeal_samples[34639]=22145;
squeal_samples[34640]=24305;
squeal_samples[34641]=26385;
squeal_samples[34642]=28355;
squeal_samples[34643]=30253;
squeal_samples[34644]=32056;
squeal_samples[34645]=33785;
squeal_samples[34646]=35425;
squeal_samples[34647]=37004;
squeal_samples[34648]=38501;
squeal_samples[34649]=39945;
squeal_samples[34650]=41311;
squeal_samples[34651]=42624;
squeal_samples[34652]=43868;
squeal_samples[34653]=45071;
squeal_samples[34654]=46209;
squeal_samples[34655]=47293;
squeal_samples[34656]=48338;
squeal_samples[34657]=49328;
squeal_samples[34658]=50284;
squeal_samples[34659]=51179;
squeal_samples[34660]=52056;
squeal_samples[34661]=52876;
squeal_samples[34662]=53671;
squeal_samples[34663]=54424;
squeal_samples[34664]=52548;
squeal_samples[34665]=46751;
squeal_samples[34666]=41262;
squeal_samples[34667]=36136;
squeal_samples[34668]=31332;
squeal_samples[34669]=26836;
squeal_samples[34670]=22630;
squeal_samples[34671]=18696;
squeal_samples[34672]=15013;
squeal_samples[34673]=11559;
squeal_samples[34674]=8337;
squeal_samples[34675]=5316;
squeal_samples[34676]=4700;
squeal_samples[34677]=7581;
squeal_samples[34678]=10392;
squeal_samples[34679]=13073;
squeal_samples[34680]=15645;
squeal_samples[34681]=18097;
squeal_samples[34682]=20439;
squeal_samples[34683]=22679;
squeal_samples[34684]=24825;
squeal_samples[34685]=26873;
squeal_samples[34686]=28833;
squeal_samples[34687]=30698;
squeal_samples[34688]=32489;
squeal_samples[34689]=34188;
squeal_samples[34690]=35819;
squeal_samples[34691]=37375;
squeal_samples[34692]=38863;
squeal_samples[34693]=40277;
squeal_samples[34694]=41634;
squeal_samples[34695]=42932;
squeal_samples[34696]=44162;
squeal_samples[34697]=45346;
squeal_samples[34698]=46476;
squeal_samples[34699]=47547;
squeal_samples[34700]=48578;
squeal_samples[34701]=49556;
squeal_samples[34702]=50499;
squeal_samples[34703]=51393;
squeal_samples[34704]=52251;
squeal_samples[34705]=53067;
squeal_samples[34706]=53851;
squeal_samples[34707]=54543;
squeal_samples[34708]=51095;
squeal_samples[34709]=45335;
squeal_samples[34710]=39939;
squeal_samples[34711]=34897;
squeal_samples[34712]=30168;
squeal_samples[34713]=25749;
squeal_samples[34714]=21605;
squeal_samples[34715]=17743;
squeal_samples[34716]=14114;
squeal_samples[34717]=10725;
squeal_samples[34718]=7553;
squeal_samples[34719]=4627;
squeal_samples[34720]=5383;
squeal_samples[34721]=8290;
squeal_samples[34722]=11058;
squeal_samples[34723]=13717;
squeal_samples[34724]=16256;
squeal_samples[34725]=18685;
squeal_samples[34726]=20996;
squeal_samples[34727]=23219;
squeal_samples[34728]=25333;
squeal_samples[34729]=27359;
squeal_samples[34730]=29295;
squeal_samples[34731]=31141;
squeal_samples[34732]=32904;
squeal_samples[34733]=34592;
squeal_samples[34734]=36204;
squeal_samples[34735]=37743;
squeal_samples[34736]=39209;
squeal_samples[34737]=40615;
squeal_samples[34738]=41954;
squeal_samples[34739]=43236;
squeal_samples[34740]=44454;
squeal_samples[34741]=45625;
squeal_samples[34742]=46733;
squeal_samples[34743]=47801;
squeal_samples[34744]=48813;
squeal_samples[34745]=49787;
squeal_samples[34746]=50715;
squeal_samples[34747]=51601;
squeal_samples[34748]=52444;
squeal_samples[34749]=53255;
squeal_samples[34750]=54030;
squeal_samples[34751]=54289;
squeal_samples[34752]=49606;
squeal_samples[34753]=43937;
squeal_samples[34754]=38638;
squeal_samples[34755]=33673;
squeal_samples[34756]=29025;
squeal_samples[34757]=24676;
squeal_samples[34758]=20603;
squeal_samples[34759]=16802;
squeal_samples[34760]=13235;
squeal_samples[34761]=9900;
squeal_samples[34762]=6779;
squeal_samples[34763]=4271;
squeal_samples[34764]=6110;
squeal_samples[34765]=8981;
squeal_samples[34766]=11726;
squeal_samples[34767]=14351;
squeal_samples[34768]=16861;
squeal_samples[34769]=19259;
squeal_samples[34770]=21552;
squeal_samples[34771]=23742;
squeal_samples[34772]=25840;
squeal_samples[34773]=27841;
squeal_samples[34774]=29751;
squeal_samples[34775]=31582;
squeal_samples[34776]=33326;
squeal_samples[34777]=34994;
squeal_samples[34778]=36583;
squeal_samples[34779]=38101;
squeal_samples[34780]=39558;
squeal_samples[34781]=40944;
squeal_samples[34782]=42271;
squeal_samples[34783]=43531;
squeal_samples[34784]=44740;
squeal_samples[34785]=45892;
squeal_samples[34786]=46998;
squeal_samples[34787]=48047;
squeal_samples[34788]=49055;
squeal_samples[34789]=50013;
squeal_samples[34790]=50928;
squeal_samples[34791]=51802;
squeal_samples[34792]=52639;
squeal_samples[34793]=53442;
squeal_samples[34794]=54203;
squeal_samples[34795]=53607;
squeal_samples[34796]=48142;
squeal_samples[34797]=42571;
squeal_samples[34798]=37353;
squeal_samples[34799]=32476;
squeal_samples[34800]=27898;
squeal_samples[34801]=23625;
squeal_samples[34802]=19619;
squeal_samples[34803]=15881;
squeal_samples[34804]=12369;
squeal_samples[34805]=9093;
squeal_samples[34806]=6016;
squeal_samples[34807]=4283;
squeal_samples[34808]=6828;
squeal_samples[34809]=9671;
squeal_samples[34810]=12383;
squeal_samples[34811]=14983;
squeal_samples[34812]=17462;
squeal_samples[34813]=19829;
squeal_samples[34814]=22101;
squeal_samples[34815]=24263;
squeal_samples[34816]=26340;
squeal_samples[34817]=28312;
squeal_samples[34818]=30209;
squeal_samples[34819]=32012;
squeal_samples[34820]=33744;
squeal_samples[34821]=35379;
squeal_samples[34822]=36962;
squeal_samples[34823]=38457;
squeal_samples[34824]=39899;
squeal_samples[34825]=41272;
squeal_samples[34826]=42577;
squeal_samples[34827]=43827;
squeal_samples[34828]=45027;
squeal_samples[34829]=46162;
squeal_samples[34830]=47254;
squeal_samples[34831]=48292;
squeal_samples[34832]=49286;
squeal_samples[34833]=50239;
squeal_samples[34834]=51136;
squeal_samples[34835]=52011;
squeal_samples[34836]=52834;
squeal_samples[34837]=53626;
squeal_samples[34838]=54378;
squeal_samples[34839]=53193;
squeal_samples[34840]=47497;
squeal_samples[34841]=41965;
squeal_samples[34842]=36786;
squeal_samples[34843]=31940;
squeal_samples[34844]=27401;
squeal_samples[34845]=23158;
squeal_samples[34846]=19178;
squeal_samples[34847]=15469;
squeal_samples[34848]=11983;
squeal_samples[34849]=8733;
squeal_samples[34850]=5681;
squeal_samples[34851]=4456;
squeal_samples[34852]=7215;
squeal_samples[34853]=10040;
squeal_samples[34854]=12736;
squeal_samples[34855]=15319;
squeal_samples[34856]=17782;
squeal_samples[34857]=20141;
squeal_samples[34858]=22391;
squeal_samples[34859]=24548;
squeal_samples[34860]=26604;
squeal_samples[34861]=28573;
squeal_samples[34862]=30453;
squeal_samples[34863]=32247;
squeal_samples[34864]=33957;
squeal_samples[34865]=35596;
squeal_samples[34866]=37158;
squeal_samples[34867]=38656;
squeal_samples[34868]=40083;
squeal_samples[34869]=41443;
squeal_samples[34870]=42749;
squeal_samples[34871]=43981;
squeal_samples[34872]=45175;
squeal_samples[34873]=46305;
squeal_samples[34874]=47387;
squeal_samples[34875]=48424;
squeal_samples[34876]=49405;
squeal_samples[34877]=50352;
squeal_samples[34878]=51253;
squeal_samples[34879]=52112;
squeal_samples[34880]=52933;
squeal_samples[34881]=53719;
squeal_samples[34882]=54472;
squeal_samples[34883]=52589;
squeal_samples[34884]=46785;
squeal_samples[34885]=41297;
squeal_samples[34886]=36164;
squeal_samples[34887]=31351;
squeal_samples[34888]=26856;
squeal_samples[34889]=22638;
squeal_samples[34890]=18703;
squeal_samples[34891]=15018;
squeal_samples[34892]=11559;
squeal_samples[34893]=8332;
squeal_samples[34894]=5306;
squeal_samples[34895]=4689;
squeal_samples[34896]=7570;
squeal_samples[34897]=10374;
squeal_samples[34898]=13061;
squeal_samples[34899]=15625;
squeal_samples[34900]=18079;
squeal_samples[34901]=20415;
squeal_samples[34902]=22657;
squeal_samples[34903]=24805;
squeal_samples[34904]=26846;
squeal_samples[34905]=28804;
squeal_samples[34906]=30668;
squeal_samples[34907]=32455;
squeal_samples[34908]=34157;
squeal_samples[34909]=35786;
squeal_samples[34910]=37343;
squeal_samples[34911]=38829;
squeal_samples[34912]=40246;
squeal_samples[34913]=41602;
squeal_samples[34914]=42894;
squeal_samples[34915]=44130;
squeal_samples[34916]=45308;
squeal_samples[34917]=46436;
squeal_samples[34918]=47513;
squeal_samples[34919]=48536;
squeal_samples[34920]=49523;
squeal_samples[34921]=50452;
squeal_samples[34922]=51352;
squeal_samples[34923]=52211;
squeal_samples[34924]=53024;
squeal_samples[34925]=53808;
squeal_samples[34926]=54552;
squeal_samples[34927]=51886;
squeal_samples[34928]=46065;
squeal_samples[34929]=40628;
squeal_samples[34930]=35527;
squeal_samples[34931]=30766;
squeal_samples[34932]=26299;
squeal_samples[34933]=22122;
squeal_samples[34934]=18224;
squeal_samples[34935]=14555;
squeal_samples[34936]=11142;
squeal_samples[34937]=7932;
squeal_samples[34938]=4938;
squeal_samples[34939]=5003;
squeal_samples[34940]=7920;
squeal_samples[34941]=10704;
squeal_samples[34942]=13378;
squeal_samples[34943]=15922;
squeal_samples[34944]=18374;
squeal_samples[34945]=20691;
squeal_samples[34946]=22925;
squeal_samples[34947]=25053;
squeal_samples[34948]=27086;
squeal_samples[34949]=29032;
squeal_samples[34950]=30885;
squeal_samples[34951]=32662;
squeal_samples[34952]=34357;
squeal_samples[34953]=35976;
squeal_samples[34954]=37523;
squeal_samples[34955]=38997;
squeal_samples[34956]=40411;
squeal_samples[34957]=41751;
squeal_samples[34958]=43043;
squeal_samples[34959]=44263;
squeal_samples[34960]=45447;
squeal_samples[34961]=46560;
squeal_samples[34962]=47633;
squeal_samples[34963]=48651;
squeal_samples[34964]=49629;
squeal_samples[34965]=50558;
squeal_samples[34966]=51450;
squeal_samples[34967]=52302;
squeal_samples[34968]=53115;
squeal_samples[34969]=53890;
squeal_samples[34970]=54587;
squeal_samples[34971]=51118;
squeal_samples[34972]=45360;
squeal_samples[34973]=39955;
squeal_samples[34974]=34908;
squeal_samples[34975]=30175;
squeal_samples[34976]=25753;
squeal_samples[34977]=21607;
squeal_samples[34978]=17738;
squeal_samples[34979]=14110;
squeal_samples[34980]=10713;
squeal_samples[34981]=7539;
squeal_samples[34982]=4609;
squeal_samples[34983]=5366;
squeal_samples[34984]=8259;
squeal_samples[34985]=11040;
squeal_samples[34986]=13689;
squeal_samples[34987]=16229;
squeal_samples[34988]=18655;
squeal_samples[34989]=20963;
squeal_samples[34990]=23188;
squeal_samples[34991]=25300;
squeal_samples[34992]=27327;
squeal_samples[34993]=29259;
squeal_samples[34994]=31103;
squeal_samples[34995]=32867;
squeal_samples[34996]=34556;
squeal_samples[34997]=36158;
squeal_samples[34998]=37704;
squeal_samples[34999]=39165;
squeal_samples[35000]=40572;
squeal_samples[35001]=41906;
squeal_samples[35002]=43187;
squeal_samples[35003]=44407;
squeal_samples[35004]=45577;
squeal_samples[35005]=46684;
squeal_samples[35006]=47754;
squeal_samples[35007]=48763;
squeal_samples[35008]=49740;
squeal_samples[35009]=50661;
squeal_samples[35010]=51548;
squeal_samples[35011]=52395;
squeal_samples[35012]=53202;
squeal_samples[35013]=53974;
squeal_samples[35014]=54503;
squeal_samples[35015]=50372;
squeal_samples[35016]=44651;
squeal_samples[35017]=39300;
squeal_samples[35018]=34288;
squeal_samples[35019]=29595;
squeal_samples[35020]=25210;
squeal_samples[35021]=21097;
squeal_samples[35022]=17262;
squeal_samples[35023]=13655;
squeal_samples[35024]=10296;
squeal_samples[35025]=7142;
squeal_samples[35026]=4380;
squeal_samples[35027]=5722;
squeal_samples[35028]=8604;
squeal_samples[35029]=11366;
squeal_samples[35030]=14003;
squeal_samples[35031]=16525;
squeal_samples[35032]=18939;
squeal_samples[35033]=21239;
squeal_samples[35034]=23440;
squeal_samples[35035]=25546;
squeal_samples[35036]=27562;
squeal_samples[35037]=29478;
squeal_samples[35038]=31325;
squeal_samples[35039]=33070;
squeal_samples[35040]=34752;
squeal_samples[35041]=36344;
squeal_samples[35042]=37876;
squeal_samples[35043]=39335;
squeal_samples[35044]=40729;
squeal_samples[35045]=42059;
squeal_samples[35046]=43333;
squeal_samples[35047]=44544;
squeal_samples[35048]=45706;
squeal_samples[35049]=46810;
squeal_samples[35050]=47872;
squeal_samples[35051]=48881;
squeal_samples[35052]=49845;
squeal_samples[35053]=50768;
squeal_samples[35054]=51643;
squeal_samples[35055]=52488;
squeal_samples[35056]=53292;
squeal_samples[35057]=54053;
squeal_samples[35058]=54316;
squeal_samples[35059]=49621;
squeal_samples[35060]=43955;
squeal_samples[35061]=38647;
squeal_samples[35062]=33670;
squeal_samples[35063]=29024;
squeal_samples[35064]=24669;
squeal_samples[35065]=20595;
squeal_samples[35066]=16788;
squeal_samples[35067]=13217;
squeal_samples[35068]=9882;
squeal_samples[35069]=6752;
squeal_samples[35070]=4239;
squeal_samples[35071]=6081;
squeal_samples[35072]=8946;
squeal_samples[35073]=11692;
squeal_samples[35074]=14315;
squeal_samples[35075]=16821;
squeal_samples[35076]=19220;
squeal_samples[35077]=21508;
squeal_samples[35078]=23701;
squeal_samples[35079]=25799;
squeal_samples[35080]=27791;
squeal_samples[35081]=29705;
squeal_samples[35082]=31533;
squeal_samples[35083]=33275;
squeal_samples[35084]=34940;
squeal_samples[35085]=36531;
squeal_samples[35086]=38047;
squeal_samples[35087]=39505;
squeal_samples[35088]=40886;
squeal_samples[35089]=42212;
squeal_samples[35090]=43475;
squeal_samples[35091]=44683;
squeal_samples[35092]=45839;
squeal_samples[35093]=46933;
squeal_samples[35094]=47995;
squeal_samples[35095]=48991;
squeal_samples[35096]=49953;
squeal_samples[35097]=50867;
squeal_samples[35098]=51744;
squeal_samples[35099]=52583;
squeal_samples[35100]=53374;
squeal_samples[35101]=54142;
squeal_samples[35102]=54017;
squeal_samples[35103]=48887;
squeal_samples[35104]=43258;
squeal_samples[35105]=37995;
squeal_samples[35106]=33064;
squeal_samples[35107]=28451;
squeal_samples[35108]=24136;
squeal_samples[35109]=20093;
squeal_samples[35110]=16317;
squeal_samples[35111]=12772;
squeal_samples[35112]=9469;
squeal_samples[35113]=6366;
squeal_samples[35114]=4198;
squeal_samples[35115]=6433;
squeal_samples[35116]=9285;
squeal_samples[35117]=12017;
squeal_samples[35118]=14624;
squeal_samples[35119]=17117;
squeal_samples[35120]=19501;
squeal_samples[35121]=21779;
squeal_samples[35122]=23958;
squeal_samples[35123]=26041;
squeal_samples[35124]=28028;
squeal_samples[35125]=29926;
squeal_samples[35126]=31746;
squeal_samples[35127]=33474;
squeal_samples[35128]=35137;
squeal_samples[35129]=36716;
squeal_samples[35130]=38226;
squeal_samples[35131]=39670;
squeal_samples[35132]=41041;
squeal_samples[35133]=42366;
squeal_samples[35134]=43620;
squeal_samples[35135]=44822;
squeal_samples[35136]=45966;
squeal_samples[35137]=47063;
squeal_samples[35138]=48104;
squeal_samples[35139]=49104;
squeal_samples[35140]=50060;
squeal_samples[35141]=50965;
squeal_samples[35142]=51839;
squeal_samples[35143]=52667;
squeal_samples[35144]=53465;
squeal_samples[35145]=54222;
squeal_samples[35146]=53617;
squeal_samples[35147]=48152;
squeal_samples[35148]=42570;
squeal_samples[35149]=37353;
squeal_samples[35150]=32463;
squeal_samples[35151]=27888;
squeal_samples[35152]=23601;
squeal_samples[35153]=19597;
squeal_samples[35154]=15846;
squeal_samples[35155]=12344;
squeal_samples[35156]=9049;
squeal_samples[35157]=5989;
squeal_samples[35158]=4233;
squeal_samples[35159]=6794;
squeal_samples[35160]=9618;
squeal_samples[35161]=12340;
squeal_samples[35162]=14933;
squeal_samples[35163]=17411;
squeal_samples[35164]=19777;
squeal_samples[35165]=22047;
squeal_samples[35166]=24212;
squeal_samples[35167]=26281;
squeal_samples[35168]=28261;
squeal_samples[35169]=30149;
squeal_samples[35170]=31952;
squeal_samples[35171]=33676;
squeal_samples[35172]=35326;
squeal_samples[35173]=36901;
squeal_samples[35174]=38395;
squeal_samples[35175]=39837;
squeal_samples[35176]=41201;
squeal_samples[35177]=42516;
squeal_samples[35178]=43762;
squeal_samples[35179]=44958;
squeal_samples[35180]=46097;
squeal_samples[35181]=47180;
squeal_samples[35182]=48228;
squeal_samples[35183]=49208;
squeal_samples[35184]=50167;
squeal_samples[35185]=51067;
squeal_samples[35186]=51936;
squeal_samples[35187]=52760;
squeal_samples[35188]=53552;
squeal_samples[35189]=54303;
squeal_samples[35190]=53696;
squeal_samples[35191]=48219;
squeal_samples[35192]=42639;
squeal_samples[35193]=37410;
squeal_samples[35194]=32518;
squeal_samples[35195]=27944;
squeal_samples[35196]=23648;
squeal_samples[35197]=19642;
squeal_samples[35198]=15890;
squeal_samples[35199]=12379;
squeal_samples[35200]=9093;
squeal_samples[35201]=6015;
squeal_samples[35202]=4267;
squeal_samples[35203]=6815;
squeal_samples[35204]=9649;
squeal_samples[35205]=12361;
squeal_samples[35206]=14956;
squeal_samples[35207]=17432;
squeal_samples[35208]=19800;
squeal_samples[35209]=22062;
squeal_samples[35210]=24230;
squeal_samples[35211]=26297;
squeal_samples[35212]=28271;
squeal_samples[35213]=30163;
squeal_samples[35214]=31966;
squeal_samples[35215]=33689;
squeal_samples[35216]=35336;
squeal_samples[35217]=36906;
squeal_samples[35218]=38408;
squeal_samples[35219]=39841;
squeal_samples[35220]=41213;
squeal_samples[35221]=42522;
squeal_samples[35222]=43768;
squeal_samples[35223]=44963;
squeal_samples[35224]=46096;
squeal_samples[35225]=47189;
squeal_samples[35226]=48225;
squeal_samples[35227]=49217;
squeal_samples[35228]=50164;
squeal_samples[35229]=51069;
squeal_samples[35230]=51937;
squeal_samples[35231]=52760;
squeal_samples[35232]=53551;
squeal_samples[35233]=54305;
squeal_samples[35234]=53694;
squeal_samples[35235]=48223;
squeal_samples[35236]=42635;
squeal_samples[35237]=37408;
squeal_samples[35238]=32511;
squeal_samples[35239]=27939;
squeal_samples[35240]=23644;
squeal_samples[35241]=19636;
squeal_samples[35242]=15885;
squeal_samples[35243]=12375;
squeal_samples[35244]=9085;
squeal_samples[35245]=6013;
squeal_samples[35246]=4259;
squeal_samples[35247]=6808;
squeal_samples[35248]=9642;
squeal_samples[35249]=12356;
squeal_samples[35250]=14945;
squeal_samples[35251]=17427;
squeal_samples[35252]=19790;
squeal_samples[35253]=22057;
squeal_samples[35254]=24225;
squeal_samples[35255]=26291;
squeal_samples[35256]=28267;
squeal_samples[35257]=30157;
squeal_samples[35258]=31956;
squeal_samples[35259]=33683;
squeal_samples[35260]=35327;
squeal_samples[35261]=36900;
squeal_samples[35262]=38398;
squeal_samples[35263]=39835;
squeal_samples[35264]=41204;
squeal_samples[35265]=42509;
squeal_samples[35266]=43759;
squeal_samples[35267]=44954;
squeal_samples[35268]=46088;
squeal_samples[35269]=47182;
squeal_samples[35270]=48209;
squeal_samples[35271]=49212;
squeal_samples[35272]=50156;
squeal_samples[35273]=51061;
squeal_samples[35274]=51924;
squeal_samples[35275]=52749;
squeal_samples[35276]=53544;
squeal_samples[35277]=54291;
squeal_samples[35278]=53687;
squeal_samples[35279]=48209;
squeal_samples[35280]=42626;
squeal_samples[35281]=37403;
squeal_samples[35282]=32501;
squeal_samples[35283]=27928;
squeal_samples[35284]=23633;
squeal_samples[35285]=19626;
squeal_samples[35286]=15874;
squeal_samples[35287]=12366;
squeal_samples[35288]=9072;
squeal_samples[35289]=6006;
squeal_samples[35290]=4245;
squeal_samples[35291]=6800;
squeal_samples[35292]=9630;
squeal_samples[35293]=12346;
squeal_samples[35294]=14934;
squeal_samples[35295]=17418;
squeal_samples[35296]=19783;
squeal_samples[35297]=22048;
squeal_samples[35298]=24214;
squeal_samples[35299]=26279;
squeal_samples[35300]=28260;
squeal_samples[35301]=30142;
squeal_samples[35302]=31950;
squeal_samples[35303]=33670;
squeal_samples[35304]=35318;
squeal_samples[35305]=36887;
squeal_samples[35306]=38391;
squeal_samples[35307]=39822;
squeal_samples[35308]=41194;
squeal_samples[35309]=42500;
squeal_samples[35310]=43746;
squeal_samples[35311]=44945;
squeal_samples[35312]=46077;
squeal_samples[35313]=47172;
squeal_samples[35314]=48198;
squeal_samples[35315]=49203;
squeal_samples[35316]=50143;
squeal_samples[35317]=51052;
squeal_samples[35318]=51913;
squeal_samples[35319]=52740;
squeal_samples[35320]=53531;
squeal_samples[35321]=54283;
squeal_samples[35322]=53674;
squeal_samples[35323]=48200;
squeal_samples[35324]=42616;
squeal_samples[35325]=37392;
squeal_samples[35326]=32490;
squeal_samples[35327]=27918;
squeal_samples[35328]=23622;
squeal_samples[35329]=19616;
squeal_samples[35330]=15864;
squeal_samples[35331]=12354;
squeal_samples[35332]=9065;
squeal_samples[35333]=5990;
squeal_samples[35334]=4240;
squeal_samples[35335]=6784;
squeal_samples[35336]=9624;
squeal_samples[35337]=12334;
squeal_samples[35338]=14924;
squeal_samples[35339]=17406;
squeal_samples[35340]=19774;
squeal_samples[35341]=22036;
squeal_samples[35342]=24205;
squeal_samples[35343]=26268;
squeal_samples[35344]=28249;
squeal_samples[35345]=30132;
squeal_samples[35346]=31939;
squeal_samples[35347]=33660;
squeal_samples[35348]=35306;
squeal_samples[35349]=36880;
squeal_samples[35350]=38376;
squeal_samples[35351]=39814;
squeal_samples[35352]=41184;
squeal_samples[35353]=42487;
squeal_samples[35354]=43739;
squeal_samples[35355]=44931;
squeal_samples[35356]=46070;
squeal_samples[35357]=47157;
squeal_samples[35358]=48193;
squeal_samples[35359]=49186;
squeal_samples[35360]=50138;
squeal_samples[35361]=51039;
squeal_samples[35362]=51903;
squeal_samples[35363]=52729;
squeal_samples[35364]=53521;
squeal_samples[35365]=54271;
squeal_samples[35366]=53666;
squeal_samples[35367]=48188;
squeal_samples[35368]=42606;
squeal_samples[35369]=37381;
squeal_samples[35370]=32480;
squeal_samples[35371]=27907;
squeal_samples[35372]=23613;
squeal_samples[35373]=19604;
squeal_samples[35374]=15854;
squeal_samples[35375]=12344;
squeal_samples[35376]=9052;
squeal_samples[35377]=5985;
squeal_samples[35378]=4223;
squeal_samples[35379]=6780;
squeal_samples[35380]=9608;
squeal_samples[35381]=12326;
squeal_samples[35382]=14914;
squeal_samples[35383]=17394;
squeal_samples[35384]=19765;
squeal_samples[35385]=22025;
squeal_samples[35386]=24193;
squeal_samples[35387]=26261;
squeal_samples[35388]=28234;
squeal_samples[35389]=30125;
squeal_samples[35390]=31927;
squeal_samples[35391]=33649;
squeal_samples[35392]=35298;
squeal_samples[35393]=36865;
squeal_samples[35394]=38369;
squeal_samples[35395]=39804;
squeal_samples[35396]=41171;
squeal_samples[35397]=42479;
squeal_samples[35398]=43727;
squeal_samples[35399]=44920;
squeal_samples[35400]=46061;
squeal_samples[35401]=47147;
squeal_samples[35402]=48180;
squeal_samples[35403]=49180;
squeal_samples[35404]=50122;
squeal_samples[35405]=51033;
squeal_samples[35406]=51889;
squeal_samples[35407]=52722;
squeal_samples[35408]=53508;
squeal_samples[35409]=54263;
squeal_samples[35410]=53653;
squeal_samples[35411]=48178;
squeal_samples[35412]=42598;
squeal_samples[35413]=37365;
squeal_samples[35414]=32478;
squeal_samples[35415]=27888;
squeal_samples[35416]=23608;
squeal_samples[35417]=19591;
squeal_samples[35418]=15844;
squeal_samples[35419]=12333;
squeal_samples[35420]=9044;
squeal_samples[35421]=5970;
squeal_samples[35422]=4217;
squeal_samples[35423]=6767;
squeal_samples[35424]=9598;
squeal_samples[35425]=12316;
squeal_samples[35426]=14902;
squeal_samples[35427]=17386;
squeal_samples[35428]=19752;
squeal_samples[35429]=22016;
squeal_samples[35430]=24183;
squeal_samples[35431]=26247;
squeal_samples[35432]=28230;
squeal_samples[35433]=30109;
squeal_samples[35434]=31918;
squeal_samples[35435]=33640;
squeal_samples[35436]=35283;
squeal_samples[35437]=36861;
squeal_samples[35438]=38354;
squeal_samples[35439]=39794;
squeal_samples[35440]=41161;
squeal_samples[35441]=42469;
squeal_samples[35442]=43714;
squeal_samples[35443]=44914;
squeal_samples[35444]=46046;
squeal_samples[35445]=47139;
squeal_samples[35446]=48169;
squeal_samples[35447]=49168;
squeal_samples[35448]=50115;
squeal_samples[35449]=51018;
squeal_samples[35450]=51883;
squeal_samples[35451]=52707;
squeal_samples[35452]=53501;
squeal_samples[35453]=54251;
squeal_samples[35454]=53642;
squeal_samples[35455]=48169;
squeal_samples[35456]=42584;
squeal_samples[35457]=37360;
squeal_samples[35458]=32460;
squeal_samples[35459]=27885;
squeal_samples[35460]=23592;
squeal_samples[35461]=19584;
squeal_samples[35462]=15831;
squeal_samples[35463]=12323;
squeal_samples[35464]=9033;
squeal_samples[35465]=5961;
squeal_samples[35466]=4206;
squeal_samples[35467]=6755;
squeal_samples[35468]=9590;
squeal_samples[35469]=12303;
squeal_samples[35470]=14893;
squeal_samples[35471]=17375;
squeal_samples[35472]=19742;
squeal_samples[35473]=22006;
squeal_samples[35474]=24170;
squeal_samples[35475]=26241;
squeal_samples[35476]=28213;
squeal_samples[35477]=30105;
squeal_samples[35478]=31903;
squeal_samples[35479]=33631;
squeal_samples[35480]=35274;
squeal_samples[35481]=36848;
squeal_samples[35482]=38345;
squeal_samples[35483]=39783;
squeal_samples[35484]=41150;
squeal_samples[35485]=42458;
squeal_samples[35486]=43706;
squeal_samples[35487]=44900;
squeal_samples[35488]=46039;
squeal_samples[35489]=47125;
squeal_samples[35490]=48162;
squeal_samples[35491]=49153;
squeal_samples[35492]=50109;
squeal_samples[35493]=51004;
squeal_samples[35494]=51874;
squeal_samples[35495]=52698;
squeal_samples[35496]=53487;
squeal_samples[35497]=54243;
squeal_samples[35498]=53630;
squeal_samples[35499]=48160;
squeal_samples[35500]=42572;
squeal_samples[35501]=37351;
squeal_samples[35502]=32448;
squeal_samples[35503]=27875;
squeal_samples[35504]=23582;
squeal_samples[35505]=19572;
squeal_samples[35506]=15822;
squeal_samples[35507]=12313;
squeal_samples[35508]=9021;
squeal_samples[35509]=5951;
squeal_samples[35510]=4195;
squeal_samples[35511]=6745;
squeal_samples[35512]=9579;
squeal_samples[35513]=12294;
squeal_samples[35514]=14880;
squeal_samples[35515]=17366;
squeal_samples[35516]=19730;
squeal_samples[35517]=21996;
squeal_samples[35518]=24161;
squeal_samples[35519]=26228;
squeal_samples[35520]=28204;
squeal_samples[35521]=30093;
squeal_samples[35522]=31894;
squeal_samples[35523]=33620;
squeal_samples[35524]=35264;
squeal_samples[35525]=36835;
squeal_samples[35526]=38338;
squeal_samples[35527]=39769;
squeal_samples[35528]=41143;
squeal_samples[35529]=42444;
squeal_samples[35530]=43698;
squeal_samples[35531]=44887;
squeal_samples[35532]=46030;
squeal_samples[35533]=47114;
squeal_samples[35534]=48150;
squeal_samples[35535]=49144;
squeal_samples[35536]=50097;
squeal_samples[35537]=50993;
squeal_samples[35538]=51865;
squeal_samples[35539]=52683;
squeal_samples[35540]=53480;
squeal_samples[35541]=54229;
squeal_samples[35542]=54099;
squeal_samples[35543]=48952;
squeal_samples[35544]=43318;
squeal_samples[35545]=38043;
squeal_samples[35546]=33105;
squeal_samples[35547]=28477;
squeal_samples[35548]=24158;
squeal_samples[35549]=20100;
squeal_samples[35550]=16320;
squeal_samples[35551]=12772;
squeal_samples[35552]=9457;
squeal_samples[35553]=6353;
squeal_samples[35554]=4168;
squeal_samples[35555]=6413;
squeal_samples[35556]=9259;
squeal_samples[35557]=11983;
squeal_samples[35558]=14589;
squeal_samples[35559]=17083;
squeal_samples[35560]=19459;
squeal_samples[35561]=21735;
squeal_samples[35562]=23911;
squeal_samples[35563]=25991;
squeal_samples[35564]=27975;
squeal_samples[35565]=29877;
squeal_samples[35566]=31687;
squeal_samples[35567]=33420;
squeal_samples[35568]=35074;
squeal_samples[35569]=36652;
squeal_samples[35570]=38162;
squeal_samples[35571]=39603;
squeal_samples[35572]=40978;
squeal_samples[35573]=42296;
squeal_samples[35574]=43548;
squeal_samples[35575]=44749;
squeal_samples[35576]=45893;
squeal_samples[35577]=46983;
squeal_samples[35578]=48028;
squeal_samples[35579]=49023;
squeal_samples[35580]=49978;
squeal_samples[35581]=50887;
squeal_samples[35582]=51758;
squeal_samples[35583]=52584;
squeal_samples[35584]=53380;
squeal_samples[35585]=54137;
squeal_samples[35586]=54381;
squeal_samples[35587]=49681;
squeal_samples[35588]=43997;
squeal_samples[35589]=38680;
squeal_samples[35590]=33701;
squeal_samples[35591]=29038;
squeal_samples[35592]=24678;
squeal_samples[35593]=20589;
squeal_samples[35594]=16778;
squeal_samples[35595]=13198;
squeal_samples[35596]=9859;
squeal_samples[35597]=6717;
squeal_samples[35598]=4205;
squeal_samples[35599]=6036;
squeal_samples[35600]=8901;
squeal_samples[35601]=11642;
squeal_samples[35602]=14262;
squeal_samples[35603]=16769;
squeal_samples[35604]=19155;
squeal_samples[35605]=21447;
squeal_samples[35606]=23636;
squeal_samples[35607]=25729;
squeal_samples[35608]=27728;
squeal_samples[35609]=29631;
squeal_samples[35610]=31455;
squeal_samples[35611]=33198;
squeal_samples[35612]=34862;
squeal_samples[35613]=36451;
squeal_samples[35614]=37968;
squeal_samples[35615]=39414;
squeal_samples[35616]=40805;
squeal_samples[35617]=42121;
squeal_samples[35618]=43387;
squeal_samples[35619]=44590;
squeal_samples[35620]=45744;
squeal_samples[35621]=46840;
squeal_samples[35622]=47893;
squeal_samples[35623]=48894;
squeal_samples[35624]=49852;
squeal_samples[35625]=50768;
squeal_samples[35626]=51638;
squeal_samples[35627]=52477;
squeal_samples[35628]=53270;
squeal_samples[35629]=54033;
squeal_samples[35630]=54551;
squeal_samples[35631]=50407;
squeal_samples[35632]=44685;
squeal_samples[35633]=39313;
squeal_samples[35634]=34299;
squeal_samples[35635]=29593;
squeal_samples[35636]=25198;
squeal_samples[35637]=21075;
squeal_samples[35638]=17231;
squeal_samples[35639]=13626;
squeal_samples[35640]=10245;
squeal_samples[35641]=7093;
squeal_samples[35642]=4319;
squeal_samples[35643]=5665;
squeal_samples[35644]=8541;
squeal_samples[35645]=11300;
squeal_samples[35646]=13932;
squeal_samples[35647]=16453;
squeal_samples[35648]=18857;
squeal_samples[35649]=21161;
squeal_samples[35650]=23358;
squeal_samples[35651]=25458;
squeal_samples[35652]=27473;
squeal_samples[35653]=29388;
squeal_samples[35654]=31221;
squeal_samples[35655]=32976;
squeal_samples[35656]=34645;
squeal_samples[35657]=36246;
squeal_samples[35658]=37773;
squeal_samples[35659]=39228;
squeal_samples[35660]=40622;
squeal_samples[35661]=41947;
squeal_samples[35662]=43220;
squeal_samples[35663]=44433;
squeal_samples[35664]=45590;
squeal_samples[35665]=46697;
squeal_samples[35666]=47750;
squeal_samples[35667]=48760;
squeal_samples[35668]=49726;
squeal_samples[35669]=50643;
squeal_samples[35670]=51527;
squeal_samples[35671]=52359;
squeal_samples[35672]=53170;
squeal_samples[35673]=53928;
squeal_samples[35674]=54616;
squeal_samples[35675]=51142;
squeal_samples[35676]=45369;
squeal_samples[35677]=39954;
squeal_samples[35678]=34897;
squeal_samples[35679]=30153;
squeal_samples[35680]=25719;
squeal_samples[35681]=21565;
squeal_samples[35682]=17686;
squeal_samples[35683]=14051;
squeal_samples[35684]=10647;
squeal_samples[35685]=7468;
squeal_samples[35686]=4528;
squeal_samples[35687]=5282;
squeal_samples[35688]=8179;
squeal_samples[35689]=10946;
squeal_samples[35690]=13595;
squeal_samples[35691]=16135;
squeal_samples[35692]=18551;
squeal_samples[35693]=20870;
squeal_samples[35694]=23074;
squeal_samples[35695]=25194;
squeal_samples[35696]=27212;
squeal_samples[35697]=29144;
squeal_samples[35698]=30989;
squeal_samples[35699]=32746;
squeal_samples[35700]=34437;
squeal_samples[35701]=36037;
squeal_samples[35702]=37579;
squeal_samples[35703]=39039;
squeal_samples[35704]=40443;
squeal_samples[35705]=41774;
squeal_samples[35706]=43055;
squeal_samples[35707]=44274;
squeal_samples[35708]=45435;
squeal_samples[35709]=46554;
squeal_samples[35710]=47612;
squeal_samples[35711]=48625;
squeal_samples[35712]=49596;
squeal_samples[35713]=50520;
squeal_samples[35714]=51405;
squeal_samples[35715]=52247;
squeal_samples[35716]=53055;
squeal_samples[35717]=53825;
squeal_samples[35718]=54567;
squeal_samples[35719]=51882;
squeal_samples[35720]=46056;
squeal_samples[35721]=40605;
squeal_samples[35722]=35496;
squeal_samples[35723]=30722;
squeal_samples[35724]=26243;
squeal_samples[35725]=22059;
squeal_samples[35726]=18150;
squeal_samples[35727]=14484;
squeal_samples[35728]=11050;
squeal_samples[35729]=7843;
squeal_samples[35730]=4837;
squeal_samples[35731]=4904;
squeal_samples[35732]=7806;
squeal_samples[35733]=10603;
squeal_samples[35734]=13254;
squeal_samples[35735]=15818;
squeal_samples[35736]=18241;
squeal_samples[35737]=20571;
squeal_samples[35738]=22793;
squeal_samples[35739]=24922;
squeal_samples[35740]=26958;
squeal_samples[35741]=28893;
squeal_samples[35742]=30753;
squeal_samples[35743]=32521;
squeal_samples[35744]=34222;
squeal_samples[35745]=35824;
squeal_samples[35746]=37381;
squeal_samples[35747]=38847;
squeal_samples[35748]=40259;
squeal_samples[35749]=41601;
squeal_samples[35750]=42888;
squeal_samples[35751]=44115;
squeal_samples[35752]=45286;
squeal_samples[35753]=46405;
squeal_samples[35754]=47472;
squeal_samples[35755]=48496;
squeal_samples[35756]=49465;
squeal_samples[35757]=50395;
squeal_samples[35758]=51286;
squeal_samples[35759]=52133;
squeal_samples[35760]=52946;
squeal_samples[35761]=53723;
squeal_samples[35762]=54468;
squeal_samples[35763]=52572;
squeal_samples[35764]=46753;
squeal_samples[35765]=41255;
squeal_samples[35766]=36108;
squeal_samples[35767]=31288;
squeal_samples[35768]=26779;
squeal_samples[35769]=22557;
squeal_samples[35770]=18612;
squeal_samples[35771]=14919;
squeal_samples[35772]=11457;
squeal_samples[35773]=8225;
squeal_samples[35774]=5189;
squeal_samples[35775]=4568;
squeal_samples[35776]=7442;
squeal_samples[35777]=10248;
squeal_samples[35778]=12922;
squeal_samples[35779]=15488;
squeal_samples[35780]=17935;
squeal_samples[35781]=20275;
squeal_samples[35782]=22514;
squeal_samples[35783]=24649;
squeal_samples[35784]=26699;
squeal_samples[35785]=28649;
squeal_samples[35786]=30513;
squeal_samples[35787]=32296;
squeal_samples[35788]=33996;
squeal_samples[35789]=35624;
squeal_samples[35790]=37173;
squeal_samples[35791]=38658;
squeal_samples[35792]=40077;
squeal_samples[35793]=41427;
squeal_samples[35794]=42723;
squeal_samples[35795]=43949;
squeal_samples[35796]=45131;
squeal_samples[35797]=46258;
squeal_samples[35798]=47331;
squeal_samples[35799]=48360;
squeal_samples[35800]=49335;
squeal_samples[35801]=50272;
squeal_samples[35802]=51164;
squeal_samples[35803]=52023;
squeal_samples[35804]=52833;
squeal_samples[35805]=53618;
squeal_samples[35806]=54361;
squeal_samples[35807]=53161;
squeal_samples[35808]=47454;
squeal_samples[35809]=41913;
squeal_samples[35810]=36720;
squeal_samples[35811]=31867;
squeal_samples[35812]=27313;
squeal_samples[35813]=23060;
squeal_samples[35814]=19077;
squeal_samples[35815]=15354;
squeal_samples[35816]=11867;
squeal_samples[35817]=8600;
squeal_samples[35818]=5550;
squeal_samples[35819]=4310;
squeal_samples[35820]=7080;
squeal_samples[35821]=9889;
squeal_samples[35822]=12588;
squeal_samples[35823]=15162;
squeal_samples[35824]=17624;
squeal_samples[35825]=19981;
squeal_samples[35826]=22225;
squeal_samples[35827]=24385;
squeal_samples[35828]=26431;
squeal_samples[35829]=28400;
squeal_samples[35830]=30271;
squeal_samples[35831]=32064;
squeal_samples[35832]=33780;
squeal_samples[35833]=35410;
squeal_samples[35834]=36975;
squeal_samples[35835]=38468;
squeal_samples[35836]=39890;
squeal_samples[35837]=41253;
squeal_samples[35838]=42550;
squeal_samples[35839]=43790;
squeal_samples[35840]=44977;
squeal_samples[35841]=46106;
squeal_samples[35842]=47187;
squeal_samples[35843]=48216;
squeal_samples[35844]=49208;
squeal_samples[35845]=50142;
squeal_samples[35846]=51049;
squeal_samples[35847]=51906;
squeal_samples[35848]=52725;
squeal_samples[35849]=53514;
squeal_samples[35850]=54255;
squeal_samples[35851]=54125;
squeal_samples[35852]=48968;
squeal_samples[35853]=43332;
squeal_samples[35854]=38044;
squeal_samples[35855]=33105;
squeal_samples[35856]=28477;
squeal_samples[35857]=24144;
squeal_samples[35858]=20094;
squeal_samples[35859]=16304;
squeal_samples[35860]=12751;
squeal_samples[35861]=9435;
squeal_samples[35862]=6323;
squeal_samples[35863]=4140;
squeal_samples[35864]=6376;
squeal_samples[35865]=9222;
squeal_samples[35866]=11947;
squeal_samples[35867]=14553;
squeal_samples[35868]=17039;
squeal_samples[35869]=19421;
squeal_samples[35870]=21689;
squeal_samples[35871]=23872;
squeal_samples[35872]=25942;
squeal_samples[35873]=27929;
squeal_samples[35874]=29829;
squeal_samples[35875]=31640;
squeal_samples[35876]=33367;
squeal_samples[35877]=35020;
squeal_samples[35878]=36602;
squeal_samples[35879]=38106;
squeal_samples[35880]=39548;
squeal_samples[35881]=40924;
squeal_samples[35882]=42237;
squeal_samples[35883]=43491;
squeal_samples[35884]=44689;
squeal_samples[35885]=45836;
squeal_samples[35886]=46925;
squeal_samples[35887]=47969;
squeal_samples[35888]=48966;
squeal_samples[35889]=49917;
squeal_samples[35890]=50825;
squeal_samples[35891]=51693;
squeal_samples[35892]=52527;
squeal_samples[35893]=53313;
squeal_samples[35894]=54076;
squeal_samples[35895]=54580;
squeal_samples[35896]=50441;
squeal_samples[35897]=44697;
squeal_samples[35898]=39333;
squeal_samples[35899]=34306;
squeal_samples[35900]=29599;
squeal_samples[35901]=25200;
squeal_samples[35902]=21076;
squeal_samples[35903]=17221;
squeal_samples[35904]=13617;
squeal_samples[35905]=10236;
squeal_samples[35906]=7076;
squeal_samples[35907]=4302;
squeal_samples[35908]=5640;
squeal_samples[35909]=8519;
squeal_samples[35910]=11272;
squeal_samples[35911]=13907;
squeal_samples[35912]=16421;
squeal_samples[35913]=18826;
squeal_samples[35914]=21129;
squeal_samples[35915]=23327;
squeal_samples[35916]=25427;
squeal_samples[35917]=27436;
squeal_samples[35918]=29350;
squeal_samples[35919]=31186;
squeal_samples[35920]=32938;
squeal_samples[35921]=34607;
squeal_samples[35922]=36207;
squeal_samples[35923]=37727;
squeal_samples[35924]=39189;
squeal_samples[35925]=40577;
squeal_samples[35926]=41907;
squeal_samples[35927]=43175;
squeal_samples[35928]=44388;
squeal_samples[35929]=45541;
squeal_samples[35930]=46649;
squeal_samples[35931]=47704;
squeal_samples[35932]=48709;
squeal_samples[35933]=49675;
squeal_samples[35934]=50590;
squeal_samples[35935]=51472;
squeal_samples[35936]=52308;
squeal_samples[35937]=53113;
squeal_samples[35938]=53879;
squeal_samples[35939]=54611;
squeal_samples[35940]=51927;
squeal_samples[35941]=46085;
squeal_samples[35942]=40634;
squeal_samples[35943]=35521;
squeal_samples[35944]=30735;
squeal_samples[35945]=26263;
squeal_samples[35946]=22071;
squeal_samples[35947]=18154;
squeal_samples[35948]=14487;
squeal_samples[35949]=11045;
squeal_samples[35950]=7837;
squeal_samples[35951]=4830;
squeal_samples[35952]=4891;
squeal_samples[35953]=7800;
squeal_samples[35954]=10582;
squeal_samples[35955]=13245;
squeal_samples[35956]=15791;
squeal_samples[35957]=18231;
squeal_samples[35958]=20546;
squeal_samples[35959]=22775;
squeal_samples[35960]=24901;
squeal_samples[35961]=26929;
squeal_samples[35962]=28871;
squeal_samples[35963]=30721;
squeal_samples[35964]=32496;
squeal_samples[35965]=34185;
squeal_samples[35966]=35803;
squeal_samples[35967]=37343;
squeal_samples[35968]=38820;
squeal_samples[35969]=40225;
squeal_samples[35970]=41570;
squeal_samples[35971]=42851;
squeal_samples[35972]=44078;
squeal_samples[35973]=45248;
squeal_samples[35974]=46367;
squeal_samples[35975]=47432;
squeal_samples[35976]=48449;
squeal_samples[35977]=49433;
squeal_samples[35978]=50354;
squeal_samples[35979]=51245;
squeal_samples[35980]=52089;
squeal_samples[35981]=52904;
squeal_samples[35982]=53679;
squeal_samples[35983]=54425;
squeal_samples[35984]=53215;
squeal_samples[35985]=47502;
squeal_samples[35986]=41953;
squeal_samples[35987]=36757;
squeal_samples[35988]=31896;
squeal_samples[35989]=27341;
squeal_samples[35990]=23082;
squeal_samples[35991]=19094;
squeal_samples[35992]=15371;
squeal_samples[35993]=11878;
squeal_samples[35994]=8608;
squeal_samples[35995]=5553;
squeal_samples[35996]=4314;
squeal_samples[35997]=7073;
squeal_samples[35998]=9885;
squeal_samples[35999]=12585;
squeal_samples[36000]=15154;
squeal_samples[36001]=17622;
squeal_samples[36002]=19969;
squeal_samples[36003]=22212;
squeal_samples[36004]=24371;
squeal_samples[36005]=26420;
squeal_samples[36006]=28387;
squeal_samples[36007]=30255;
squeal_samples[36008]=32052;
squeal_samples[36009]=33753;
squeal_samples[36010]=35401;
squeal_samples[36011]=36949;
squeal_samples[36012]=38449;
squeal_samples[36013]=39865;
squeal_samples[36014]=41229;
squeal_samples[36015]=42527;
squeal_samples[36016]=43765;
squeal_samples[36017]=44953;
squeal_samples[36018]=46080;
squeal_samples[36019]=47159;
squeal_samples[36020]=48192;
squeal_samples[36021]=49178;
squeal_samples[36022]=50119;
squeal_samples[36023]=51016;
squeal_samples[36024]=51873;
squeal_samples[36025]=52696;
squeal_samples[36026]=53478;
squeal_samples[36027]=54229;
squeal_samples[36028]=54088;
squeal_samples[36029]=48940;
squeal_samples[36030]=43291;
squeal_samples[36031]=38017;
squeal_samples[36032]=33068;
squeal_samples[36033]=28444;
squeal_samples[36034]=24109;
squeal_samples[36035]=20059;
squeal_samples[36036]=16265;
squeal_samples[36037]=12715;
squeal_samples[36038]=9396;
squeal_samples[36039]=6288;
squeal_samples[36040]=4102;
squeal_samples[36041]=6337;
squeal_samples[36042]=9188;
squeal_samples[36043]=11906;
squeal_samples[36044]=14520;
squeal_samples[36045]=16998;
squeal_samples[36046]=19386;
squeal_samples[36047]=21652;
squeal_samples[36048]=23828;
squeal_samples[36049]=25906;
squeal_samples[36050]=27890;
squeal_samples[36051]=29789;
squeal_samples[36052]=31596;
squeal_samples[36053]=33329;
squeal_samples[36054]=34985;
squeal_samples[36055]=36561;
squeal_samples[36056]=38068;
squeal_samples[36057]=39508;
squeal_samples[36058]=40881;
squeal_samples[36059]=42196;
squeal_samples[36060]=43447;
squeal_samples[36061]=44647;
squeal_samples[36062]=45794;
squeal_samples[36063]=46881;
squeal_samples[36064]=47927;
squeal_samples[36065]=48923;
squeal_samples[36066]=49876;
squeal_samples[36067]=50780;
squeal_samples[36068]=51653;
squeal_samples[36069]=52481;
squeal_samples[36070]=53274;
squeal_samples[36071]=54031;
squeal_samples[36072]=54545;
squeal_samples[36073]=50396;
squeal_samples[36074]=44661;
squeal_samples[36075]=39291;
squeal_samples[36076]=34267;
squeal_samples[36077]=29559;
squeal_samples[36078]=25155;
squeal_samples[36079]=21035;
squeal_samples[36080]=17177;
squeal_samples[36081]=13574;
squeal_samples[36082]=10195;
squeal_samples[36083]=7032;
squeal_samples[36084]=4261;
squeal_samples[36085]=5597;
squeal_samples[36086]=8475;
squeal_samples[36087]=11231;
squeal_samples[36088]=13862;
squeal_samples[36089]=16382;
squeal_samples[36090]=18781;
squeal_samples[36091]=21088;
squeal_samples[36092]=23283;
squeal_samples[36093]=25385;
squeal_samples[36094]=27393;
squeal_samples[36095]=29308;
squeal_samples[36096]=31143;
squeal_samples[36097]=32896;
squeal_samples[36098]=34565;
squeal_samples[36099]=36163;
squeal_samples[36100]=37684;
squeal_samples[36101]=39148;
squeal_samples[36102]=40533;
squeal_samples[36103]=41866;
squeal_samples[36104]=43131;
squeal_samples[36105]=44346;
squeal_samples[36106]=45497;
squeal_samples[36107]=46609;
squeal_samples[36108]=47658;
squeal_samples[36109]=48670;
squeal_samples[36110]=49629;
squeal_samples[36111]=50550;
squeal_samples[36112]=51427;
squeal_samples[36113]=52267;
squeal_samples[36114]=53071;
squeal_samples[36115]=53834;
squeal_samples[36116]=54572;
squeal_samples[36117]=51880;
squeal_samples[36118]=46046;
squeal_samples[36119]=40591;
squeal_samples[36120]=35476;
squeal_samples[36121]=30695;
squeal_samples[36122]=26220;
squeal_samples[36123]=22027;
squeal_samples[36124]=18114;
squeal_samples[36125]=14442;
squeal_samples[36126]=11004;
squeal_samples[36127]=7794;
squeal_samples[36128]=4787;
squeal_samples[36129]=4848;
squeal_samples[36130]=7758;
squeal_samples[36131]=10539;
squeal_samples[36132]=13204;
squeal_samples[36133]=15746;
squeal_samples[36134]=18190;
squeal_samples[36135]=20503;
squeal_samples[36136]=22731;
squeal_samples[36137]=24861;
squeal_samples[36138]=26885;
squeal_samples[36139]=28828;
squeal_samples[36140]=30680;
squeal_samples[36141]=32452;
squeal_samples[36142]=34143;
squeal_samples[36143]=35760;
squeal_samples[36144]=37301;
squeal_samples[36145]=38778;
squeal_samples[36146]=40180;
squeal_samples[36147]=41532;
squeal_samples[36148]=42803;
squeal_samples[36149]=44040;
squeal_samples[36150]=45203;
squeal_samples[36151]=46325;
squeal_samples[36152]=47389;
squeal_samples[36153]=48409;
squeal_samples[36154]=49386;
squeal_samples[36155]=50315;
squeal_samples[36156]=51200;
squeal_samples[36157]=52049;
squeal_samples[36158]=52860;
squeal_samples[36159]=53637;
squeal_samples[36160]=54381;
squeal_samples[36161]=53173;
squeal_samples[36162]=47461;
squeal_samples[36163]=41909;
squeal_samples[36164]=36715;
squeal_samples[36165]=31852;
squeal_samples[36166]=27300;
squeal_samples[36167]=23038;
squeal_samples[36168]=19054;
squeal_samples[36169]=15324;
squeal_samples[36170]=11840;
squeal_samples[36171]=8561;
squeal_samples[36172]=5515;
squeal_samples[36173]=4268;
squeal_samples[36174]=7031;
squeal_samples[36175]=9845;
squeal_samples[36176]=12539;
squeal_samples[36177]=15114;
squeal_samples[36178]=17578;
squeal_samples[36179]=19926;
squeal_samples[36180]=22171;
squeal_samples[36181]=24328;
squeal_samples[36182]=26377;
squeal_samples[36183]=28343;
squeal_samples[36184]=30216;
squeal_samples[36185]=32005;
squeal_samples[36186]=33715;
squeal_samples[36187]=35353;
squeal_samples[36188]=36912;
squeal_samples[36189]=38401;
squeal_samples[36190]=39826;
squeal_samples[36191]=41185;
squeal_samples[36192]=42483;
squeal_samples[36193]=43726;
squeal_samples[36194]=44908;
squeal_samples[36195]=46036;
squeal_samples[36196]=47119;
squeal_samples[36197]=48147;
squeal_samples[36198]=49136;
squeal_samples[36199]=50078;
squeal_samples[36200]=50970;
squeal_samples[36201]=51833;
squeal_samples[36202]=52651;
squeal_samples[36203]=53436;
squeal_samples[36204]=54184;
squeal_samples[36205]=54422;
squeal_samples[36206]=49710;
squeal_samples[36207]=44018;
squeal_samples[36208]=38681;
squeal_samples[36209]=33693;
squeal_samples[36210]=29020;
squeal_samples[36211]=24653;
squeal_samples[36212]=20560;
squeal_samples[36213]=16737;
squeal_samples[36214]=13152;
squeal_samples[36215]=9801;
squeal_samples[36216]=6663;
squeal_samples[36217]=4134;
squeal_samples[36218]=5971;
squeal_samples[36219]=8826;
squeal_samples[36220]=11570;
squeal_samples[36221]=14183;
squeal_samples[36222]=16690;
squeal_samples[36223]=19071;
squeal_samples[36224]=21365;
squeal_samples[36225]=23545;
squeal_samples[36226]=25634;
squeal_samples[36227]=27633;
squeal_samples[36228]=29537;
squeal_samples[36229]=31353;
squeal_samples[36230]=33100;
squeal_samples[36231]=34753;
squeal_samples[36232]=36351;
squeal_samples[36233]=37856;
squeal_samples[36234]=39312;
squeal_samples[36235]=40685;
squeal_samples[36236]=42013;
squeal_samples[36237]=43268;
squeal_samples[36238]=44476;
squeal_samples[36239]=45623;
squeal_samples[36240]=46723;
squeal_samples[36241]=47767;
squeal_samples[36242]=48773;
squeal_samples[36243]=49730;
squeal_samples[36244]=50640;
squeal_samples[36245]=51516;
squeal_samples[36246]=52349;
squeal_samples[36247]=53140;
squeal_samples[36248]=53908;
squeal_samples[36249]=54636;
squeal_samples[36250]=51941;
squeal_samples[36251]=46100;
squeal_samples[36252]=40641;
squeal_samples[36253]=35519;
squeal_samples[36254]=30741;
squeal_samples[36255]=26250;
squeal_samples[36256]=22057;
squeal_samples[36257]=18135;
squeal_samples[36258]=14464;
squeal_samples[36259]=11027;
squeal_samples[36260]=7810;
squeal_samples[36261]=4799;
squeal_samples[36262]=4859;
squeal_samples[36263]=7765;
squeal_samples[36264]=10543;
squeal_samples[36265]=13211;
squeal_samples[36266]=15752;
squeal_samples[36267]=18190;
squeal_samples[36268]=20505;
squeal_samples[36269]=22730;
squeal_samples[36270]=24856;
squeal_samples[36271]=26881;
squeal_samples[36272]=28824;
squeal_samples[36273]=30674;
squeal_samples[36274]=32447;
squeal_samples[36275]=34133;
squeal_samples[36276]=35749;
squeal_samples[36277]=37293;
squeal_samples[36278]=38759;
squeal_samples[36279]=40174;
squeal_samples[36280]=41511;
squeal_samples[36281]=42798;
squeal_samples[36282]=44018;
squeal_samples[36283]=45192;
squeal_samples[36284]=46308;
squeal_samples[36285]=47373;
squeal_samples[36286]=48394;
squeal_samples[36287]=49362;
squeal_samples[36288]=50297;
squeal_samples[36289]=51182;
squeal_samples[36290]=52034;
squeal_samples[36291]=52838;
squeal_samples[36292]=53616;
squeal_samples[36293]=54353;
squeal_samples[36294]=53735;
squeal_samples[36295]=48235;
squeal_samples[36296]=42641;
squeal_samples[36297]=37387;
squeal_samples[36298]=32483;
squeal_samples[36299]=27888;
squeal_samples[36300]=23585;
squeal_samples[36301]=19566;
squeal_samples[36302]=15799;
squeal_samples[36303]=12276;
squeal_samples[36304]=8980;
squeal_samples[36305]=5897;
squeal_samples[36306]=4134;
squeal_samples[36307]=6686;
squeal_samples[36308]=9504;
squeal_samples[36309]=12218;
squeal_samples[36310]=14801;
squeal_samples[36311]=17279;
squeal_samples[36312]=19635;
squeal_samples[36313]=21903;
squeal_samples[36314]=24061;
squeal_samples[36315]=26122;
squeal_samples[36316]=28097;
squeal_samples[36317]=29979;
squeal_samples[36318]=31782;
squeal_samples[36319]=33496;
squeal_samples[36320]=35145;
squeal_samples[36321]=36708;
squeal_samples[36322]=38211;
squeal_samples[36323]=39638;
squeal_samples[36324]=41010;
squeal_samples[36325]=42308;
squeal_samples[36326]=43559;
squeal_samples[36327]=44746;
squeal_samples[36328]=45885;
squeal_samples[36329]=46973;
squeal_samples[36330]=48006;
squeal_samples[36331]=48997;
squeal_samples[36332]=49941;
squeal_samples[36333]=50842;
squeal_samples[36334]=51707;
squeal_samples[36335]=52528;
squeal_samples[36336]=53317;
squeal_samples[36337]=54070;
squeal_samples[36338]=54580;
squeal_samples[36339]=50423;
squeal_samples[36340]=44680;
squeal_samples[36341]=39307;
squeal_samples[36342]=34276;
squeal_samples[36343]=29562;
squeal_samples[36344]=25160;
squeal_samples[36345]=21027;
squeal_samples[36346]=17177;
squeal_samples[36347]=13562;
squeal_samples[36348]=10181;
squeal_samples[36349]=7016;
squeal_samples[36350]=4241;
squeal_samples[36351]=5577;
squeal_samples[36352]=8455;
squeal_samples[36353]=11204;
squeal_samples[36354]=13833;
squeal_samples[36355]=16353;
squeal_samples[36356]=18752;
squeal_samples[36357]=21056;
squeal_samples[36358]=23246;
squeal_samples[36359]=25350;
squeal_samples[36360]=27355;
squeal_samples[36361]=29271;
squeal_samples[36362]=31108;
squeal_samples[36363]=32851;
squeal_samples[36364]=34526;
squeal_samples[36365]=36120;
squeal_samples[36366]=37641;
squeal_samples[36367]=39103;
squeal_samples[36368]=40487;
squeal_samples[36369]=41821;
squeal_samples[36370]=43084;
squeal_samples[36371]=44297;
squeal_samples[36372]=45452;
squeal_samples[36373]=46558;
squeal_samples[36374]=47613;
squeal_samples[36375]=48616;
squeal_samples[36376]=49583;
squeal_samples[36377]=50500;
squeal_samples[36378]=51377;
squeal_samples[36379]=52212;
squeal_samples[36380]=53018;
squeal_samples[36381]=53781;
squeal_samples[36382]=54512;
squeal_samples[36383]=52616;
squeal_samples[36384]=46782;
squeal_samples[36385]=41268;
squeal_samples[36386]=36116;
squeal_samples[36387]=31286;
squeal_samples[36388]=26766;
squeal_samples[36389]=22533;
squeal_samples[36390]=18582;
squeal_samples[36391]=14877;
squeal_samples[36392]=11414;
squeal_samples[36393]=8170;
squeal_samples[36394]=5132;
squeal_samples[36395]=4500;
squeal_samples[36396]=7379;
squeal_samples[36397]=10178;
squeal_samples[36398]=12849;
squeal_samples[36399]=15415;
squeal_samples[36400]=17857;
squeal_samples[36401]=20191;
squeal_samples[36402]=22430;
squeal_samples[36403]=24559;
squeal_samples[36404]=26604;
squeal_samples[36405]=28555;
squeal_samples[36406]=30418;
squeal_samples[36407]=32197;
squeal_samples[36408]=33893;
squeal_samples[36409]=35521;
squeal_samples[36410]=37066;
squeal_samples[36411]=38554;
squeal_samples[36412]=39964;
squeal_samples[36413]=41319;
squeal_samples[36414]=42607;
squeal_samples[36415]=43844;
squeal_samples[36416]=45009;
squeal_samples[36417]=46140;
squeal_samples[36418]=47207;
squeal_samples[36419]=48239;
squeal_samples[36420]=49212;
squeal_samples[36421]=50149;
squeal_samples[36422]=51045;
squeal_samples[36423]=51891;
squeal_samples[36424]=52709;
squeal_samples[36425]=53486;
squeal_samples[36426]=54234;
squeal_samples[36427]=54094;
squeal_samples[36428]=48933;
squeal_samples[36429]=43285;
squeal_samples[36430]=38000;
squeal_samples[36431]=33047;
squeal_samples[36432]=28415;
squeal_samples[36433]=24081;
squeal_samples[36434]=20022;
squeal_samples[36435]=16229;
squeal_samples[36436]=12677;
squeal_samples[36437]=9345;
squeal_samples[36438]=6239;
squeal_samples[36439]=4047;
squeal_samples[36440]=6288;
squeal_samples[36441]=9128;
squeal_samples[36442]=11851;
squeal_samples[36443]=14454;
squeal_samples[36444]=16943;
squeal_samples[36445]=19321;
squeal_samples[36446]=21590;
squeal_samples[36447]=23765;
squeal_samples[36448]=25838;
squeal_samples[36449]=27821;
squeal_samples[36450]=29720;
squeal_samples[36451]=31528;
squeal_samples[36452]=33258;
squeal_samples[36453]=34907;
squeal_samples[36454]=36492;
squeal_samples[36455]=37990;
squeal_samples[36456]=39437;
squeal_samples[36457]=40806;
squeal_samples[36458]=42124;
squeal_samples[36459]=43370;
squeal_samples[36460]=44574;
squeal_samples[36461]=45707;
squeal_samples[36462]=46809;
squeal_samples[36463]=47842;
squeal_samples[36464]=48848;
squeal_samples[36465]=49793;
squeal_samples[36466]=50705;
squeal_samples[36467]=51564;
squeal_samples[36468]=52400;
squeal_samples[36469]=53186;
squeal_samples[36470]=53946;
squeal_samples[36471]=54619;
squeal_samples[36472]=51135;
squeal_samples[36473]=45350;
squeal_samples[36474]=39928;
squeal_samples[36475]=34855;
squeal_samples[36476]=30105;
squeal_samples[36477]=25662;
squeal_samples[36478]=21503;
squeal_samples[36479]=17617;
squeal_samples[36480]=13970;
squeal_samples[36481]=10563;
squeal_samples[36482]=7370;
squeal_samples[36483]=4432;
squeal_samples[36484]=5176;
squeal_samples[36485]=8070;
squeal_samples[36486]=10835;
squeal_samples[36487]=13481;
squeal_samples[36488]=16012;
squeal_samples[36489]=18433;
squeal_samples[36490]=20742;
squeal_samples[36491]=22949;
squeal_samples[36492]=25061;
squeal_samples[36493]=27081;
squeal_samples[36494]=29007;
squeal_samples[36495]=30845;
squeal_samples[36496]=32613;
squeal_samples[36497]=34282;
squeal_samples[36498]=35897;
squeal_samples[36499]=37425;
squeal_samples[36500]=38895;
squeal_samples[36501]=40285;
squeal_samples[36502]=41625;
squeal_samples[36503]=42894;
squeal_samples[36504]=44122;
squeal_samples[36505]=45274;
squeal_samples[36506]=46397;
squeal_samples[36507]=47446;
squeal_samples[36508]=48467;
squeal_samples[36509]=49432;
squeal_samples[36510]=50353;
squeal_samples[36511]=51238;
squeal_samples[36512]=52079;
squeal_samples[36513]=52892;
squeal_samples[36514]=53653;
squeal_samples[36515]=54395;
squeal_samples[36516]=53761;
squeal_samples[36517]=48265;
squeal_samples[36518]=42664;
squeal_samples[36519]=37404;
squeal_samples[36520]=32503;
squeal_samples[36521]=27896;
squeal_samples[36522]=23597;
squeal_samples[36523]=19563;
squeal_samples[36524]=15804;
squeal_samples[36525]=12271;
squeal_samples[36526]=8970;
squeal_samples[36527]=5882;
squeal_samples[36528]=4123;
squeal_samples[36529]=6659;
squeal_samples[36530]=9497;
squeal_samples[36531]=12191;
squeal_samples[36532]=14787;
squeal_samples[36533]=17254;
squeal_samples[36534]=19619;
squeal_samples[36535]=21873;
squeal_samples[36536]=24038;
squeal_samples[36537]=26097;
squeal_samples[36538]=28069;
squeal_samples[36539]=29953;
squeal_samples[36540]=31750;
squeal_samples[36541]=33469;
squeal_samples[36542]=35111;
squeal_samples[36543]=36680;
squeal_samples[36544]=38177;
squeal_samples[36545]=39605;
squeal_samples[36546]=40969;
squeal_samples[36547]=42276;
squeal_samples[36548]=43519;
squeal_samples[36549]=44712;
squeal_samples[36550]=45842;
squeal_samples[36551]=46930;
squeal_samples[36552]=47967;
squeal_samples[36553]=48953;
squeal_samples[36554]=49899;
squeal_samples[36555]=50802;
squeal_samples[36556]=51663;
squeal_samples[36557]=52487;
squeal_samples[36558]=53275;
squeal_samples[36559]=54026;
squeal_samples[36560]=54697;
squeal_samples[36561]=51206;
squeal_samples[36562]=45416;
squeal_samples[36563]=39987;
squeal_samples[36564]=34913;
squeal_samples[36565]=30151;
squeal_samples[36566]=25708;
squeal_samples[36567]=21542;
squeal_samples[36568]=17647;
squeal_samples[36569]=14003;
squeal_samples[36570]=10585;
squeal_samples[36571]=7398;
squeal_samples[36572]=4449;
squeal_samples[36573]=5198;
squeal_samples[36574]=8082;
squeal_samples[36575]=10856;
squeal_samples[36576]=13495;
squeal_samples[36577]=16032;
squeal_samples[36578]=18442;
squeal_samples[36579]=20755;
squeal_samples[36580]=22953;
squeal_samples[36581]=25070;
squeal_samples[36582]=27086;
squeal_samples[36583]=29012;
squeal_samples[36584]=30854;
squeal_samples[36585]=32609;
squeal_samples[36586]=34294;
squeal_samples[36587]=35892;
squeal_samples[36588]=37431;
squeal_samples[36589]=38885;
squeal_samples[36590]=40292;
squeal_samples[36591]=41618;
squeal_samples[36592]=42902;
squeal_samples[36593]=44111;
squeal_samples[36594]=45275;
squeal_samples[36595]=46388;
squeal_samples[36596]=47443;
squeal_samples[36597]=48457;
squeal_samples[36598]=49421;
squeal_samples[36599]=50345;
squeal_samples[36600]=51229;
squeal_samples[36601]=52075;
squeal_samples[36602]=52875;
squeal_samples[36603]=53650;
squeal_samples[36604]=54379;
squeal_samples[36605]=53754;
squeal_samples[36606]=48250;
squeal_samples[36607]=42645;
squeal_samples[36608]=37399;
squeal_samples[36609]=32482;
squeal_samples[36610]=27885;
squeal_samples[36611]=23579;
squeal_samples[36612]=19549;
squeal_samples[36613]=15787;
squeal_samples[36614]=12257;
squeal_samples[36615]=8953;
squeal_samples[36616]=5868;
squeal_samples[36617]=4106;
squeal_samples[36618]=6645;
squeal_samples[36619]=9475;
squeal_samples[36620]=12176;
squeal_samples[36621]=14765;
squeal_samples[36622]=17240;
squeal_samples[36623]=19596;
squeal_samples[36624]=21855;
squeal_samples[36625]=24015;
squeal_samples[36626]=26076;
squeal_samples[36627]=28050;
squeal_samples[36628]=29928;
squeal_samples[36629]=31735;
squeal_samples[36630]=33449;
squeal_samples[36631]=35093;
squeal_samples[36632]=36656;
squeal_samples[36633]=38160;
squeal_samples[36634]=39585;
squeal_samples[36635]=40954;
squeal_samples[36636]=42254;
squeal_samples[36637]=43504;
squeal_samples[36638]=44687;
squeal_samples[36639]=45829;
squeal_samples[36640]=46909;
squeal_samples[36641]=47944;
squeal_samples[36642]=48935;
squeal_samples[36643]=49876;
squeal_samples[36644]=50787;
squeal_samples[36645]=51642;
squeal_samples[36646]=52473;
squeal_samples[36647]=53252;
squeal_samples[36648]=54008;
squeal_samples[36649]=54672;
squeal_samples[36650]=51188;
squeal_samples[36651]=45394;
squeal_samples[36652]=39966;
squeal_samples[36653]=34893;
squeal_samples[36654]=30134;
squeal_samples[36655]=25689;
squeal_samples[36656]=21519;
squeal_samples[36657]=17629;
squeal_samples[36658]=13984;
squeal_samples[36659]=10567;
squeal_samples[36660]=7376;
squeal_samples[36661]=4429;
squeal_samples[36662]=5181;
squeal_samples[36663]=8064;
squeal_samples[36664]=10831;
squeal_samples[36665]=13480;
squeal_samples[36666]=16005;
squeal_samples[36667]=18426;
squeal_samples[36668]=20731;
squeal_samples[36669]=22940;
squeal_samples[36670]=25048;
squeal_samples[36671]=27064;
squeal_samples[36672]=28994;
squeal_samples[36673]=30830;
squeal_samples[36674]=32591;
squeal_samples[36675]=34271;
squeal_samples[36676]=35874;
squeal_samples[36677]=37406;
squeal_samples[36678]=38869;
squeal_samples[36679]=40266;
squeal_samples[36680]=41603;
squeal_samples[36681]=42877;
squeal_samples[36682]=44092;
squeal_samples[36683]=45254;
squeal_samples[36684]=46366;
squeal_samples[36685]=47424;
squeal_samples[36686]=48435;
squeal_samples[36687]=49400;
squeal_samples[36688]=50324;
squeal_samples[36689]=51210;
squeal_samples[36690]=52051;
squeal_samples[36691]=52857;
squeal_samples[36692]=53626;
squeal_samples[36693]=54362;
squeal_samples[36694]=53729;
squeal_samples[36695]=48234;
squeal_samples[36696]=42619;
squeal_samples[36697]=37383;
squeal_samples[36698]=32458;
squeal_samples[36699]=27867;
squeal_samples[36700]=23555;
squeal_samples[36701]=19531;
squeal_samples[36702]=15765;
squeal_samples[36703]=12235;
squeal_samples[36704]=8935;
squeal_samples[36705]=5845;
squeal_samples[36706]=4086;
squeal_samples[36707]=6626;
squeal_samples[36708]=9450;
squeal_samples[36709]=12159;
squeal_samples[36710]=14743;
squeal_samples[36711]=17219;
squeal_samples[36712]=19576;
squeal_samples[36713]=21833;
squeal_samples[36714]=23996;
squeal_samples[36715]=26054;
squeal_samples[36716]=28030;
squeal_samples[36717]=29912;
squeal_samples[36718]=31713;
squeal_samples[36719]=33431;
squeal_samples[36720]=35070;
squeal_samples[36721]=36638;
squeal_samples[36722]=38136;
squeal_samples[36723]=39566;
squeal_samples[36724]=40932;
squeal_samples[36725]=42235;
squeal_samples[36726]=43482;
squeal_samples[36727]=44667;
squeal_samples[36728]=45807;
squeal_samples[36729]=46889;
squeal_samples[36730]=47923;
squeal_samples[36731]=48914;
squeal_samples[36732]=49856;
squeal_samples[36733]=50765;
squeal_samples[36734]=51623;
squeal_samples[36735]=52450;
squeal_samples[36736]=53232;
squeal_samples[36737]=53988;
squeal_samples[36738]=54650;
squeal_samples[36739]=51170;
squeal_samples[36740]=45370;
squeal_samples[36741]=39948;
squeal_samples[36742]=34870;
squeal_samples[36743]=30114;
squeal_samples[36744]=25669;
squeal_samples[36745]=21497;
squeal_samples[36746]=17610;
squeal_samples[36747]=13961;
squeal_samples[36748]=10549;
squeal_samples[36749]=7351;
squeal_samples[36750]=4413;
squeal_samples[36751]=5156;
squeal_samples[36752]=8047;
squeal_samples[36753]=10808;
squeal_samples[36754]=13459;
squeal_samples[36755]=15986;
squeal_samples[36756]=18404;
squeal_samples[36757]=20710;
squeal_samples[36758]=22920;
squeal_samples[36759]=25026;
squeal_samples[36760]=27046;
squeal_samples[36761]=28970;
squeal_samples[36762]=30813;
squeal_samples[36763]=32566;
squeal_samples[36764]=34255;
squeal_samples[36765]=35848;
squeal_samples[36766]=37390;
squeal_samples[36767]=38845;
squeal_samples[36768]=40248;
squeal_samples[36769]=41580;
squeal_samples[36770]=42858;
squeal_samples[36771]=44069;
squeal_samples[36772]=45235;
squeal_samples[36773]=46345;
squeal_samples[36774]=47403;
squeal_samples[36775]=48416;
squeal_samples[36776]=49377;
squeal_samples[36777]=50305;
squeal_samples[36778]=51188;
squeal_samples[36779]=52032;
squeal_samples[36780]=52836;
squeal_samples[36781]=53605;
squeal_samples[36782]=54341;
squeal_samples[36783]=53710;
squeal_samples[36784]=48210;
squeal_samples[36785]=42603;
squeal_samples[36786]=37358;
squeal_samples[36787]=32439;
squeal_samples[36788]=27846;
squeal_samples[36789]=23535;
squeal_samples[36790]=19509;
squeal_samples[36791]=15746;
squeal_samples[36792]=12213;
squeal_samples[36793]=8914;
squeal_samples[36794]=5826;
squeal_samples[36795]=4063;
squeal_samples[36796]=6606;
squeal_samples[36797]=9430;
squeal_samples[36798]=12138;
squeal_samples[36799]=14722;
squeal_samples[36800]=17199;
squeal_samples[36801]=19554;
squeal_samples[36802]=21814;
squeal_samples[36803]=23973;
squeal_samples[36804]=26037;
squeal_samples[36805]=28004;
squeal_samples[36806]=29897;
squeal_samples[36807]=31688;
squeal_samples[36808]=33414;
squeal_samples[36809]=35046;
squeal_samples[36810]=36619;
squeal_samples[36811]=38114;
squeal_samples[36812]=39547;
squeal_samples[36813]=40911;
squeal_samples[36814]=42214;
squeal_samples[36815]=43461;
squeal_samples[36816]=44647;
squeal_samples[36817]=45785;
squeal_samples[36818]=46871;
squeal_samples[36819]=47899;
squeal_samples[36820]=48896;
squeal_samples[36821]=49834;
squeal_samples[36822]=50745;
squeal_samples[36823]=51602;
squeal_samples[36824]=52429;
squeal_samples[36825]=53212;
squeal_samples[36826]=53966;
squeal_samples[36827]=54632;
squeal_samples[36828]=51146;
squeal_samples[36829]=45351;
squeal_samples[36830]=39927;
squeal_samples[36831]=34848;
squeal_samples[36832]=30097;
squeal_samples[36833]=25644;
squeal_samples[36834]=21479;
squeal_samples[36835]=17587;
squeal_samples[36836]=13943;
squeal_samples[36837]=10526;
squeal_samples[36838]=7332;
squeal_samples[36839]=4391;
squeal_samples[36840]=5136;
squeal_samples[36841]=8025;
squeal_samples[36842]=10789;
squeal_samples[36843]=13438;
squeal_samples[36844]=15964;
squeal_samples[36845]=18385;
squeal_samples[36846]=20688;
squeal_samples[36847]=22900;
squeal_samples[36848]=25006;
squeal_samples[36849]=27024;
squeal_samples[36850]=28950;
squeal_samples[36851]=30792;
squeal_samples[36852]=32546;
squeal_samples[36853]=34233;
squeal_samples[36854]=35829;
squeal_samples[36855]=37367;
squeal_samples[36856]=38828;
squeal_samples[36857]=40222;
squeal_samples[36858]=41565;
squeal_samples[36859]=42831;
squeal_samples[36860]=44054;
squeal_samples[36861]=45211;
squeal_samples[36862]=46325;
squeal_samples[36863]=47384;
squeal_samples[36864]=48390;
squeal_samples[36865]=49363;
squeal_samples[36866]=50278;
squeal_samples[36867]=51172;
squeal_samples[36868]=52006;
squeal_samples[36869]=52820;
squeal_samples[36870]=53580;
squeal_samples[36871]=54322;
squeal_samples[36872]=54166;
squeal_samples[36873]=48998;
squeal_samples[36874]=43339;
squeal_samples[36875]=38040;
squeal_samples[36876]=33086;
squeal_samples[36877]=28438;
squeal_samples[36878]=24101;
squeal_samples[36879]=20027;
squeal_samples[36880]=16231;
squeal_samples[36881]=12672;
squeal_samples[36882]=9337;
squeal_samples[36883]=6224;
squeal_samples[36884]=4027;
squeal_samples[36885]=6257;
squeal_samples[36886]=9101;
squeal_samples[36887]=11819;
squeal_samples[36888]=14416;
squeal_samples[36889]=16910;
squeal_samples[36890]=19270;
squeal_samples[36891]=21551;
squeal_samples[36892]=23712;
squeal_samples[36893]=25789;
squeal_samples[36894]=27772;
squeal_samples[36895]=29664;
squeal_samples[36896]=31472;
squeal_samples[36897]=33203;
squeal_samples[36898]=34847;
squeal_samples[36899]=36425;
squeal_samples[36900]=37929;
squeal_samples[36901]=39371;
squeal_samples[36902]=40740;
squeal_samples[36903]=42051;
squeal_samples[36904]=43302;
squeal_samples[36905]=44495;
squeal_samples[36906]=45644;
squeal_samples[36907]=46723;
squeal_samples[36908]=47773;
squeal_samples[36909]=48759;
squeal_samples[36910]=49715;
squeal_samples[36911]=50618;
squeal_samples[36912]=51489;
squeal_samples[36913]=52316;
squeal_samples[36914]=53104;
squeal_samples[36915]=53862;
squeal_samples[36916]=54588;
squeal_samples[36917]=52674;
squeal_samples[36918]=46831;
squeal_samples[36919]=41306;
squeal_samples[36920]=36142;
squeal_samples[36921]=31302;
squeal_samples[36922]=26777;
squeal_samples[36923]=22531;
squeal_samples[36924]=18573;
squeal_samples[36925]=14858;
squeal_samples[36926]=11395;
squeal_samples[36927]=8134;
squeal_samples[36928]=5100;
squeal_samples[36929]=4457;
squeal_samples[36930]=7335;
squeal_samples[36931]=10128;
squeal_samples[36932]=12802;
squeal_samples[36933]=15358;
squeal_samples[36934]=17804;
squeal_samples[36935]=20130;
squeal_samples[36936]=22365;
squeal_samples[36937]=24494;
squeal_samples[36938]=26539;
squeal_samples[36939]=28483;
squeal_samples[36940]=30348;
squeal_samples[36941]=32119;
squeal_samples[36942]=33821;
squeal_samples[36943]=35440;
squeal_samples[36944]=36989;
squeal_samples[36945]=38467;
squeal_samples[36946]=39882;
squeal_samples[36947]=41229;
squeal_samples[36948]=42517;
squeal_samples[36949]=43748;
squeal_samples[36950]=44920;
squeal_samples[36951]=46043;
squeal_samples[36952]=47120;
squeal_samples[36953]=48136;
squeal_samples[36954]=49117;
squeal_samples[36955]=50051;
squeal_samples[36956]=50937;
squeal_samples[36957]=51799;
squeal_samples[36958]=52599;
squeal_samples[36959]=53387;
squeal_samples[36960]=54128;
squeal_samples[36961]=54623;
squeal_samples[36962]=50464;
squeal_samples[36963]=44704;
squeal_samples[36964]=39323;
squeal_samples[36965]=34276;
squeal_samples[36966]=29563;
squeal_samples[36967]=25140;
squeal_samples[36968]=21009;
squeal_samples[36969]=17142;
squeal_samples[36970]=13526;
squeal_samples[36971]=10137;
squeal_samples[36972]=6964;
squeal_samples[36973]=4182;
squeal_samples[36974]=5510;
squeal_samples[36975]=8388;
squeal_samples[36976]=11131;
squeal_samples[36977]=13764;
squeal_samples[36978]=16279;
squeal_samples[36979]=18669;
squeal_samples[36980]=20972;
squeal_samples[36981]=23164;
squeal_samples[36982]=25263;
squeal_samples[36983]=27264;
squeal_samples[36984]=29180;
squeal_samples[36985]=31010;
squeal_samples[36986]=32755;
squeal_samples[36987]=34428;
squeal_samples[36988]=36017;
squeal_samples[36989]=37541;
squeal_samples[36990]=38997;
squeal_samples[36991]=40382;
squeal_samples[36992]=41712;
squeal_samples[36993]=42970;
squeal_samples[36994]=44185;
squeal_samples[36995]=45337;
squeal_samples[36996]=46440;
squeal_samples[36997]=47494;
squeal_samples[36998]=48502;
squeal_samples[36999]=49466;
squeal_samples[37000]=50373;
squeal_samples[37001]=51260;
squeal_samples[37002]=52090;
squeal_samples[37003]=52896;
squeal_samples[37004]=53654;
squeal_samples[37005]=54388;
squeal_samples[37006]=53751;
squeal_samples[37007]=48249;
squeal_samples[37008]=42634;
squeal_samples[37009]=37380;
squeal_samples[37010]=32461;
squeal_samples[37011]=27862;
squeal_samples[37012]=23549;
squeal_samples[37013]=19518;
squeal_samples[37014]=15746;
squeal_samples[37015]=12220;
squeal_samples[37016]=8907;
squeal_samples[37017]=5820;
squeal_samples[37018]=4052;
squeal_samples[37019]=6601;
squeal_samples[37020]=9420;
squeal_samples[37021]=12125;
squeal_samples[37022]=14708;
squeal_samples[37023]=17179;
squeal_samples[37024]=19536;
squeal_samples[37025]=21794;
squeal_samples[37026]=23955;
squeal_samples[37027]=26016;
squeal_samples[37028]=27988;
squeal_samples[37029]=29863;
squeal_samples[37030]=31667;
squeal_samples[37031]=33380;
squeal_samples[37032]=35021;
squeal_samples[37033]=36585;
squeal_samples[37034]=38087;
squeal_samples[37035]=39509;
squeal_samples[37036]=40882;
squeal_samples[37037]=42179;
squeal_samples[37038]=43425;
squeal_samples[37039]=44611;
squeal_samples[37040]=45747;
squeal_samples[37041]=46831;
squeal_samples[37042]=47869;
squeal_samples[37043]=48856;
squeal_samples[37044]=49800;
squeal_samples[37045]=50704;
squeal_samples[37046]=51561;
squeal_samples[37047]=52388;
squeal_samples[37048]=53172;
squeal_samples[37049]=53922;
squeal_samples[37050]=54646;
squeal_samples[37051]=51942;
squeal_samples[37052]=46088;
squeal_samples[37053]=40613;
squeal_samples[37054]=35486;
squeal_samples[37055]=30691;
squeal_samples[37056]=26202;
squeal_samples[37057]=21996;
squeal_samples[37058]=18068;
squeal_samples[37059]=14386;
squeal_samples[37060]=10939;
squeal_samples[37061]=7725;
squeal_samples[37062]=4699;
squeal_samples[37063]=4755;
squeal_samples[37064]=7658;
squeal_samples[37065]=10438;
squeal_samples[37066]=13097;
squeal_samples[37067]=15638;
squeal_samples[37068]=18070;
squeal_samples[37069]=20384;
squeal_samples[37070]=22604;
squeal_samples[37071]=24723;
squeal_samples[37072]=26759;
squeal_samples[37073]=28684;
squeal_samples[37074]=30541;
squeal_samples[37075]=32305;
squeal_samples[37076]=33995;
squeal_samples[37077]=35607;
squeal_samples[37078]=37145;
squeal_samples[37079]=38618;
squeal_samples[37080]=40022;
squeal_samples[37081]=41362;
squeal_samples[37082]=42645;
squeal_samples[37083]=43867;
squeal_samples[37084]=45037;
squeal_samples[37085]=46148;
squeal_samples[37086]=47217;
squeal_samples[37087]=48234;
squeal_samples[37088]=49202;
squeal_samples[37089]=50135;
squeal_samples[37090]=51018;
squeal_samples[37091]=51866;
squeal_samples[37092]=52677;
squeal_samples[37093]=53450;
squeal_samples[37094]=54186;
squeal_samples[37095]=54415;
squeal_samples[37096]=49691;
squeal_samples[37097]=43981;
squeal_samples[37098]=38642;
squeal_samples[37099]=33641;
squeal_samples[37100]=28960;
squeal_samples[37101]=24576;
squeal_samples[37102]=20480;
squeal_samples[37103]=16649;
squeal_samples[37104]=13056;
squeal_samples[37105]=9699;
squeal_samples[37106]=6552;
squeal_samples[37107]=4019;
squeal_samples[37108]=5846;
squeal_samples[37109]=8709;
squeal_samples[37110]=11438;
squeal_samples[37111]=14054;
squeal_samples[37112]=16550;
squeal_samples[37113]=18934;
squeal_samples[37114]=21221;
squeal_samples[37115]=23400;
squeal_samples[37116]=25488;
squeal_samples[37117]=27476;
squeal_samples[37118]=29385;
squeal_samples[37119]=31199;
squeal_samples[37120]=32937;
squeal_samples[37121]=34597;
squeal_samples[37122]=36182;
squeal_samples[37123]=37696;
squeal_samples[37124]=39138;
squeal_samples[37125]=40521;
squeal_samples[37126]=41842;
squeal_samples[37127]=43098;
squeal_samples[37128]=44300;
squeal_samples[37129]=45447;
squeal_samples[37130]=46546;
squeal_samples[37131]=47592;
squeal_samples[37132]=48592;
squeal_samples[37133]=49547;
squeal_samples[37134]=50458;
squeal_samples[37135]=51330;
squeal_samples[37136]=52161;
squeal_samples[37137]=52959;
squeal_samples[37138]=53719;
squeal_samples[37139]=54442;
squeal_samples[37140]=53227;
squeal_samples[37141]=47496;
squeal_samples[37142]=41930;
squeal_samples[37143]=36717;
squeal_samples[37144]=31841;
squeal_samples[37145]=27269;
squeal_samples[37146]=23001;
squeal_samples[37147]=19000;
squeal_samples[37148]=15261;
squeal_samples[37149]=11758;
squeal_samples[37150]=8482;
squeal_samples[37151]=5418;
squeal_samples[37152]=4170;
squeal_samples[37153]=6926;
squeal_samples[37154]=9734;
squeal_samples[37155]=12424;
squeal_samples[37156]=14992;
squeal_samples[37157]=17454;
squeal_samples[37158]=19791;
squeal_samples[37159]=22042;
squeal_samples[37160]=24182;
squeal_samples[37161]=26237;
squeal_samples[37162]=28194;
squeal_samples[37163]=30067;
squeal_samples[37164]=31854;
squeal_samples[37165]=33558;
squeal_samples[37166]=35193;
squeal_samples[37167]=36742;
squeal_samples[37168]=38237;
squeal_samples[37169]=39652;
squeal_samples[37170]=41013;
squeal_samples[37171]=42305;
squeal_samples[37172]=43547;
squeal_samples[37173]=44726;
squeal_samples[37174]=45857;
squeal_samples[37175]=46932;
squeal_samples[37176]=47960;
squeal_samples[37177]=48946;
squeal_samples[37178]=49884;
squeal_samples[37179]=50780;
squeal_samples[37180]=51641;
squeal_samples[37181]=52453;
squeal_samples[37182]=53239;
squeal_samples[37183]=53986;
squeal_samples[37184]=54648;
squeal_samples[37185]=51154;
squeal_samples[37186]=45353;
squeal_samples[37187]=39922;
squeal_samples[37188]=34845;
squeal_samples[37189]=30077;
squeal_samples[37190]=25628;
squeal_samples[37191]=21457;
squeal_samples[37192]=17562;
squeal_samples[37193]=13910;
squeal_samples[37194]=10492;
squeal_samples[37195]=7299;
squeal_samples[37196]=4352;
squeal_samples[37197]=5091;
squeal_samples[37198]=7986;
squeal_samples[37199]=10745;
squeal_samples[37200]=13391;
squeal_samples[37201]=15917;
squeal_samples[37202]=18332;
squeal_samples[37203]=20641;
squeal_samples[37204]=22843;
squeal_samples[37205]=24957;
squeal_samples[37206]=26966;
squeal_samples[37207]=28898;
squeal_samples[37208]=30733;
squeal_samples[37209]=32494;
squeal_samples[37210]=34169;
squeal_samples[37211]=35771;
squeal_samples[37212]=37304;
squeal_samples[37213]=38767;
squeal_samples[37214]=40158;
squeal_samples[37215]=41495;
squeal_samples[37216]=42769;
squeal_samples[37217]=43984;
squeal_samples[37218]=45146;
squeal_samples[37219]=46254;
squeal_samples[37220]=47315;
squeal_samples[37221]=48328;
squeal_samples[37222]=49291;
squeal_samples[37223]=50217;
squeal_samples[37224]=51096;
squeal_samples[37225]=51938;
squeal_samples[37226]=52744;
squeal_samples[37227]=53511;
squeal_samples[37228]=54247;
squeal_samples[37229]=54471;
squeal_samples[37230]=49736;
squeal_samples[37231]=44025;
squeal_samples[37232]=38685;
squeal_samples[37233]=33669;
squeal_samples[37234]=29000;
squeal_samples[37235]=24600;
squeal_samples[37236]=20507;
squeal_samples[37237]=16664;
squeal_samples[37238]=13076;
squeal_samples[37239]=9709;
squeal_samples[37240]=6566;
squeal_samples[37241]=4025;
squeal_samples[37242]=5854;
squeal_samples[37243]=8710;
squeal_samples[37244]=11439;
squeal_samples[37245]=14058;
squeal_samples[37246]=16547;
squeal_samples[37247]=18941;
squeal_samples[37248]=21212;
squeal_samples[37249]=23401;
squeal_samples[37250]=25481;
squeal_samples[37251]=27474;
squeal_samples[37252]=29373;
squeal_samples[37253]=31192;
squeal_samples[37254]=32927;
squeal_samples[37255]=34588;
squeal_samples[37256]=36173;
squeal_samples[37257]=37684;
squeal_samples[37258]=39131;
squeal_samples[37259]=40506;
squeal_samples[37260]=41826;
squeal_samples[37261]=43085;
squeal_samples[37262]=44282;
squeal_samples[37263]=45436;
squeal_samples[37264]=46528;
squeal_samples[37265]=47573;
squeal_samples[37266]=48572;
squeal_samples[37267]=49526;
squeal_samples[37268]=50438;
squeal_samples[37269]=51311;
squeal_samples[37270]=52136;
squeal_samples[37271]=52939;
squeal_samples[37272]=53694;
squeal_samples[37273]=54423;
squeal_samples[37274]=53789;
squeal_samples[37275]=48271;
squeal_samples[37276]=42657;
squeal_samples[37277]=37390;
squeal_samples[37278]=32479;
squeal_samples[37279]=27862;
squeal_samples[37280]=23550;
squeal_samples[37281]=19513;
squeal_samples[37282]=15739;
squeal_samples[37283]=12206;
squeal_samples[37284]=8896;
squeal_samples[37285]=5804;
squeal_samples[37286]=4039;
squeal_samples[37287]=6570;
squeal_samples[37288]=9401;
squeal_samples[37289]=12099;
squeal_samples[37290]=14679;
squeal_samples[37291]=17151;
squeal_samples[37292]=19505;
squeal_samples[37293]=21766;
squeal_samples[37294]=23918;
squeal_samples[37295]=25984;
squeal_samples[37296]=27945;
squeal_samples[37297]=29831;
squeal_samples[37298]=31625;
squeal_samples[37299]=33341;
squeal_samples[37300]=34978;
squeal_samples[37301]=36549;
squeal_samples[37302]=38043;
squeal_samples[37303]=39472;
squeal_samples[37304]=40833;
squeal_samples[37305]=42135;
squeal_samples[37306]=43380;
squeal_samples[37307]=44563;
squeal_samples[37308]=45705;
squeal_samples[37309]=46781;
squeal_samples[37310]=47820;
squeal_samples[37311]=48804;
squeal_samples[37312]=49750;
squeal_samples[37313]=50652;
squeal_samples[37314]=51510;
squeal_samples[37315]=52335;
squeal_samples[37316]=53122;
squeal_samples[37317]=53870;
squeal_samples[37318]=54596;
squeal_samples[37319]=52670;
squeal_samples[37320]=46826;
squeal_samples[37321]=41296;
squeal_samples[37322]=36122;
squeal_samples[37323]=31284;
squeal_samples[37324]=26744;
squeal_samples[37325]=22508;
squeal_samples[37326]=18537;
squeal_samples[37327]=14821;
squeal_samples[37328]=11349;
squeal_samples[37329]=8091;
squeal_samples[37330]=5051;
squeal_samples[37331]=4408;
squeal_samples[37332]=7278;
squeal_samples[37333]=10075;
squeal_samples[37334]=12745;
squeal_samples[37335]=15300;
squeal_samples[37336]=17742;
squeal_samples[37337]=20071;
squeal_samples[37338]=22303;
squeal_samples[37339]=24435;
squeal_samples[37340]=26473;
squeal_samples[37341]=28417;
squeal_samples[37342]=30277;
squeal_samples[37343]=32053;
squeal_samples[37344]=33750;
squeal_samples[37345]=35368;
squeal_samples[37346]=36920;
squeal_samples[37347]=38393;
squeal_samples[37348]=39813;
squeal_samples[37349]=41151;
squeal_samples[37350]=42440;
squeal_samples[37351]=43673;
squeal_samples[37352]=44841;
squeal_samples[37353]=45970;
squeal_samples[37354]=47033;
squeal_samples[37355]=48065;
squeal_samples[37356]=49036;
squeal_samples[37357]=49969;
squeal_samples[37358]=50859;
squeal_samples[37359]=51710;
squeal_samples[37360]=52524;
squeal_samples[37361]=53299;
squeal_samples[37362]=54048;
squeal_samples[37363]=54704;
squeal_samples[37364]=51205;
squeal_samples[37365]=45397;
squeal_samples[37366]=39960;
squeal_samples[37367]=34870;
squeal_samples[37368]=30109;
squeal_samples[37369]=25650;
squeal_samples[37370]=21481;
squeal_samples[37371]=17577;
squeal_samples[37372]=13921;
squeal_samples[37373]=10505;
squeal_samples[37374]=7307;
squeal_samples[37375]=4353;
squeal_samples[37376]=5094;
squeal_samples[37377]=7982;
squeal_samples[37378]=10742;
squeal_samples[37379]=13382;
squeal_samples[37380]=15909;
squeal_samples[37381]=18322;
squeal_samples[37382]=20627;
squeal_samples[37383]=22834;
squeal_samples[37384]=24943;
squeal_samples[37385]=26953;
squeal_samples[37386]=28881;
squeal_samples[37387]=30722;
squeal_samples[37388]=32472;
squeal_samples[37389]=34151;
squeal_samples[37390]=35750;
squeal_samples[37391]=37280;
squeal_samples[37392]=38747;
squeal_samples[37393]=40139;
squeal_samples[37394]=41475;
squeal_samples[37395]=42743;
squeal_samples[37396]=43962;
squeal_samples[37397]=45117;
squeal_samples[37398]=46232;
squeal_samples[37399]=47283;
squeal_samples[37400]=48302;
squeal_samples[37401]=49264;
squeal_samples[37402]=50182;
squeal_samples[37403]=51069;
squeal_samples[37404]=51905;
squeal_samples[37405]=52715;
squeal_samples[37406]=53478;
squeal_samples[37407]=54221;
squeal_samples[37408]=54430;
squeal_samples[37409]=49709;
squeal_samples[37410]=43993;
squeal_samples[37411]=38648;
squeal_samples[37412]=33642;
squeal_samples[37413]=28961;
squeal_samples[37414]=24566;
squeal_samples[37415]=20469;
squeal_samples[37416]=16630;
squeal_samples[37417]=13039;
squeal_samples[37418]=9674;
squeal_samples[37419]=6530;
squeal_samples[37420]=3988;
squeal_samples[37421]=5820;
squeal_samples[37422]=8671;
squeal_samples[37423]=11407;
squeal_samples[37424]=14018;
squeal_samples[37425]=16515;
squeal_samples[37426]=18897;
squeal_samples[37427]=21177;
squeal_samples[37428]=23365;
squeal_samples[37429]=25444;
squeal_samples[37430]=27434;
squeal_samples[37431]=29338;
squeal_samples[37432]=31154;
squeal_samples[37433]=32892;
squeal_samples[37434]=34546;
squeal_samples[37435]=36132;
squeal_samples[37436]=37644;
squeal_samples[37437]=39088;
squeal_samples[37438]=40465;
squeal_samples[37439]=41786;
squeal_samples[37440]=43041;
squeal_samples[37441]=44251;
squeal_samples[37442]=45388;
squeal_samples[37443]=46493;
squeal_samples[37444]=47534;
squeal_samples[37445]=48536;
squeal_samples[37446]=49491;
squeal_samples[37447]=50397;
squeal_samples[37448]=51274;
squeal_samples[37449]=52102;
squeal_samples[37450]=52901;
squeal_samples[37451]=53653;
squeal_samples[37452]=54385;
squeal_samples[37453]=53742;
squeal_samples[37454]=48235;
squeal_samples[37455]=42617;
squeal_samples[37456]=37353;
squeal_samples[37457]=32434;
squeal_samples[37458]=27824;
squeal_samples[37459]=23510;
squeal_samples[37460]=19475;
squeal_samples[37461]=15697;
squeal_samples[37462]=12164;
squeal_samples[37463]=8855;
squeal_samples[37464]=5763;
squeal_samples[37465]=3996;
squeal_samples[37466]=6531;
squeal_samples[37467]=9358;
squeal_samples[37468]=12057;
squeal_samples[37469]=14644;
squeal_samples[37470]=17110;
squeal_samples[37471]=19463;
squeal_samples[37472]=21725;
squeal_samples[37473]=23877;
squeal_samples[37474]=25941;
squeal_samples[37475]=27912;
squeal_samples[37476]=29787;
squeal_samples[37477]=31585;
squeal_samples[37478]=33299;
squeal_samples[37479]=34942;
squeal_samples[37480]=36508;
squeal_samples[37481]=38001;
squeal_samples[37482]=39432;
squeal_samples[37483]=40790;
squeal_samples[37484]=42095;
squeal_samples[37485]=43336;
squeal_samples[37486]=44525;
squeal_samples[37487]=45661;
squeal_samples[37488]=46741;
squeal_samples[37489]=47779;
squeal_samples[37490]=48760;
squeal_samples[37491]=49712;
squeal_samples[37492]=50608;
squeal_samples[37493]=51475;
squeal_samples[37494]=52294;
squeal_samples[37495]=53080;
squeal_samples[37496]=53830;
squeal_samples[37497]=54552;
squeal_samples[37498]=52632;
squeal_samples[37499]=46782;
squeal_samples[37500]=41257;
squeal_samples[37501]=36079;
squeal_samples[37502]=31243;
squeal_samples[37503]=26704;
squeal_samples[37504]=22464;
squeal_samples[37505]=18497;
squeal_samples[37506]=14780;
squeal_samples[37507]=11306;
squeal_samples[37508]=8052;
squeal_samples[37509]=5008;
squeal_samples[37510]=4365;
squeal_samples[37511]=7240;
squeal_samples[37512]=10031;
squeal_samples[37513]=12705;
squeal_samples[37514]=15259;
squeal_samples[37515]=17699;
squeal_samples[37516]=20032;
squeal_samples[37517]=22260;
squeal_samples[37518]=24395;
squeal_samples[37519]=26429;
squeal_samples[37520]=28379;
squeal_samples[37521]=30232;
squeal_samples[37522]=32015;
squeal_samples[37523]=33706;
squeal_samples[37524]=35329;
squeal_samples[37525]=36875;
squeal_samples[37526]=38357;
squeal_samples[37527]=39764;
squeal_samples[37528]=41117;
squeal_samples[37529]=42394;
squeal_samples[37530]=43634;
squeal_samples[37531]=44798;
squeal_samples[37532]=45928;
squeal_samples[37533]=46994;
squeal_samples[37534]=48020;
squeal_samples[37535]=48998;
squeal_samples[37536]=49924;
squeal_samples[37537]=50819;
squeal_samples[37538]=51669;
squeal_samples[37539]=52481;
squeal_samples[37540]=53257;
squeal_samples[37541]=54006;
squeal_samples[37542]=54715;
squeal_samples[37543]=52003;
squeal_samples[37544]=46136;
squeal_samples[37545]=40651;
squeal_samples[37546]=35519;
squeal_samples[37547]=30708;
squeal_samples[37548]=26210;
squeal_samples[37549]=22002;
squeal_samples[37550]=18057;
squeal_samples[37551]=14378;
squeal_samples[37552]=10918;
squeal_samples[37553]=7694;
squeal_samples[37554]=4672;
squeal_samples[37555]=4719;
squeal_samples[37556]=7621;
squeal_samples[37557]=10394;
squeal_samples[37558]=13056;
squeal_samples[37559]=15586;
squeal_samples[37560]=18019;
squeal_samples[37561]=20332;
squeal_samples[37562]=22551;
squeal_samples[37563]=24665;
squeal_samples[37564]=26691;
squeal_samples[37565]=28627;
squeal_samples[37566]=30475;
squeal_samples[37567]=32233;
squeal_samples[37568]=33927;
squeal_samples[37569]=35533;
squeal_samples[37570]=37072;
squeal_samples[37571]=38542;
squeal_samples[37572]=39944;
squeal_samples[37573]=41289;
squeal_samples[37574]=42559;
squeal_samples[37575]=43784;
squeal_samples[37576]=44949;
squeal_samples[37577]=46066;
squeal_samples[37578]=47131;
squeal_samples[37579]=48145;
squeal_samples[37580]=49118;
squeal_samples[37581]=50040;
squeal_samples[37582]=50926;
squeal_samples[37583]=51774;
squeal_samples[37584]=52583;
squeal_samples[37585]=53352;
squeal_samples[37586]=54093;
squeal_samples[37587]=54744;
squeal_samples[37588]=51241;
squeal_samples[37589]=45431;
squeal_samples[37590]=39989;
squeal_samples[37591]=34895;
squeal_samples[37592]=30126;
squeal_samples[37593]=25666;
squeal_samples[37594]=21485;
squeal_samples[37595]=17587;
squeal_samples[37596]=13922;
squeal_samples[37597]=10504;
squeal_samples[37598]=7296;
squeal_samples[37599]=4346;
squeal_samples[37600]=5080;
squeal_samples[37601]=7966;
squeal_samples[37602]=10732;
squeal_samples[37603]=13364;
squeal_samples[37604]=15896;
squeal_samples[37605]=18304;
squeal_samples[37606]=20607;
squeal_samples[37607]=22810;
squeal_samples[37608]=24916;
squeal_samples[37609]=26930;
squeal_samples[37610]=28855;
squeal_samples[37611]=30694;
squeal_samples[37612]=32444;
squeal_samples[37613]=34123;
squeal_samples[37614]=35718;
squeal_samples[37615]=37251;
squeal_samples[37616]=38711;
squeal_samples[37617]=40102;
squeal_samples[37618]=41440;
squeal_samples[37619]=42708;
squeal_samples[37620]=43924;
squeal_samples[37621]=45086;
squeal_samples[37622]=46190;
squeal_samples[37623]=47253;
squeal_samples[37624]=48257;
squeal_samples[37625]=49230;
squeal_samples[37626]=50141;
squeal_samples[37627]=51027;
squeal_samples[37628]=51864;
squeal_samples[37629]=52674;
squeal_samples[37630]=53436;
squeal_samples[37631]=54173;
squeal_samples[37632]=54656;
squeal_samples[37633]=50488;
squeal_samples[37634]=44718;
squeal_samples[37635]=39323;
squeal_samples[37636]=34269;
squeal_samples[37637]=29543;
squeal_samples[37638]=25114;
squeal_samples[37639]=20974;
squeal_samples[37640]=17101;
squeal_samples[37641]=13473;
squeal_samples[37642]=10082;
squeal_samples[37643]=6896;
squeal_samples[37644]=4118;
squeal_samples[37645]=5434;
squeal_samples[37646]=8315;
squeal_samples[37647]=11051;
squeal_samples[37648]=13680;
squeal_samples[37649]=16193;
squeal_samples[37650]=18582;
squeal_samples[37651]=20877;
squeal_samples[37652]=23072;
squeal_samples[37653]=25166;
squeal_samples[37654]=27164;
squeal_samples[37655]=29079;
squeal_samples[37656]=30902;
squeal_samples[37657]=32650;
squeal_samples[37658]=34316;
squeal_samples[37659]=35905;
squeal_samples[37660]=37430;
squeal_samples[37661]=38878;
squeal_samples[37662]=40268;
squeal_samples[37663]=41590;
squeal_samples[37664]=42858;
squeal_samples[37665]=44057;
squeal_samples[37666]=45218;
squeal_samples[37667]=46316;
squeal_samples[37668]=47370;
squeal_samples[37669]=48377;
squeal_samples[37670]=49326;
squeal_samples[37671]=50252;
squeal_samples[37672]=51118;
squeal_samples[37673]=51963;
squeal_samples[37674]=52757;
squeal_samples[37675]=53522;
squeal_samples[37676]=54253;
squeal_samples[37677]=54468;
squeal_samples[37678]=49731;
squeal_samples[37679]=44015;
squeal_samples[37680]=38663;
squeal_samples[37681]=33655;
squeal_samples[37682]=28958;
squeal_samples[37683]=24575;
squeal_samples[37684]=20461;
squeal_samples[37685]=16626;
squeal_samples[37686]=13027;
squeal_samples[37687]=9663;
squeal_samples[37688]=6510;
squeal_samples[37689]=3969;
squeal_samples[37690]=5796;
squeal_samples[37691]=8646;
squeal_samples[37692]=11382;
squeal_samples[37693]=13989;
squeal_samples[37694]=16485;
squeal_samples[37695]=18866;
squeal_samples[37696]=21144;
squeal_samples[37697]=23327;
squeal_samples[37698]=25412;
squeal_samples[37699]=27395;
squeal_samples[37700]=29305;
squeal_samples[37701]=31113;
squeal_samples[37702]=32850;
squeal_samples[37703]=34508;
squeal_samples[37704]=36088;
squeal_samples[37705]=37606;
squeal_samples[37706]=39046;
squeal_samples[37707]=40424;
squeal_samples[37708]=41745;
squeal_samples[37709]=42995;
squeal_samples[37710]=44204;
squeal_samples[37711]=45345;
squeal_samples[37712]=46443;
squeal_samples[37713]=47485;
squeal_samples[37714]=48483;
squeal_samples[37715]=49439;
squeal_samples[37716]=50353;
squeal_samples[37717]=51219;
squeal_samples[37718]=52054;
squeal_samples[37719]=52845;
squeal_samples[37720]=53605;
squeal_samples[37721]=54328;
squeal_samples[37722]=54173;
squeal_samples[37723]=48984;
squeal_samples[37724]=43316;
squeal_samples[37725]=38007;
squeal_samples[37726]=33040;
squeal_samples[37727]=28384;
squeal_samples[37728]=24038;
squeal_samples[37729]=19956;
squeal_samples[37730]=16155;
squeal_samples[37731]=12581;
squeal_samples[37732]=9246;
squeal_samples[37733]=6119;
squeal_samples[37734]=3920;
squeal_samples[37735]=6152;
squeal_samples[37736]=8981;
squeal_samples[37737]=11705;
squeal_samples[37738]=14298;
squeal_samples[37739]=16779;
squeal_samples[37740]=19149;
squeal_samples[37741]=21416;
squeal_samples[37742]=23582;
squeal_samples[37743]=25656;
squeal_samples[37744]=27632;
squeal_samples[37745]=29519;
squeal_samples[37746]=31327;
squeal_samples[37747]=33051;
squeal_samples[37748]=34703;
squeal_samples[37749]=36275;
squeal_samples[37750]=37777;
squeal_samples[37751]=39211;
squeal_samples[37752]=40582;
squeal_samples[37753]=41891;
squeal_samples[37754]=43139;
squeal_samples[37755]=44338;
squeal_samples[37756]=45474;
squeal_samples[37757]=46567;
squeal_samples[37758]=47601;
squeal_samples[37759]=48600;
squeal_samples[37760]=49542;
squeal_samples[37761]=50450;
squeal_samples[37762]=51312;
squeal_samples[37763]=52143;
squeal_samples[37764]=52926;
squeal_samples[37765]=53686;
squeal_samples[37766]=54408;
squeal_samples[37767]=53762;
squeal_samples[37768]=48250;
squeal_samples[37769]=42624;
squeal_samples[37770]=37356;
squeal_samples[37771]=32432;
squeal_samples[37772]=27815;
squeal_samples[37773]=23500;
squeal_samples[37774]=19459;
squeal_samples[37775]=15679;
squeal_samples[37776]=12146;
squeal_samples[37777]=8830;
squeal_samples[37778]=5735;
squeal_samples[37779]=3965;
squeal_samples[37780]=6503;
squeal_samples[37781]=9321;
squeal_samples[37782]=12025;
squeal_samples[37783]=14602;
squeal_samples[37784]=17074;
squeal_samples[37785]=19425;
squeal_samples[37786]=21683;
squeal_samples[37787]=23838;
squeal_samples[37788]=25895;
squeal_samples[37789]=27865;
squeal_samples[37790]=29743;
squeal_samples[37791]=31538;
squeal_samples[37792]=33255;
squeal_samples[37793]=34889;
squeal_samples[37794]=36458;
squeal_samples[37795]=37944;
squeal_samples[37796]=39375;
squeal_samples[37797]=40739;
squeal_samples[37798]=42039;
squeal_samples[37799]=43284;
squeal_samples[37800]=44470;
squeal_samples[37801]=45600;
squeal_samples[37802]=46690;
squeal_samples[37803]=47717;
squeal_samples[37804]=48709;
squeal_samples[37805]=49650;
squeal_samples[37806]=50548;
squeal_samples[37807]=51413;
squeal_samples[37808]=52231;
squeal_samples[37809]=53019;
squeal_samples[37810]=53765;
squeal_samples[37811]=54486;
squeal_samples[37812]=53253;
squeal_samples[37813]=47515;
squeal_samples[37814]=41936;
squeal_samples[37815]=36714;
squeal_samples[37816]=31833;
squeal_samples[37817]=27247;
squeal_samples[37818]=22971;
squeal_samples[37819]=18958;
squeal_samples[37820]=15220;
squeal_samples[37821]=11704;
squeal_samples[37822]=8426;
squeal_samples[37823]=5345;
squeal_samples[37824]=4101;
squeal_samples[37825]=6847;
squeal_samples[37826]=9658;
squeal_samples[37827]=12336;
squeal_samples[37828]=14909;
squeal_samples[37829]=17362;
squeal_samples[37830]=19701;
squeal_samples[37831]=21945;
squeal_samples[37832]=24088;
squeal_samples[37833]=26133;
squeal_samples[37834]=28096;
squeal_samples[37835]=29957;
squeal_samples[37836]=31748;
squeal_samples[37837]=33446;
squeal_samples[37838]=35080;
squeal_samples[37839]=36631;
squeal_samples[37840]=38124;
squeal_samples[37841]=39533;
squeal_samples[37842]=40896;
squeal_samples[37843]=42188;
squeal_samples[37844]=43423;
squeal_samples[37845]=44603;
squeal_samples[37846]=45734;
squeal_samples[37847]=46807;
squeal_samples[37848]=47834;
squeal_samples[37849]=48816;
squeal_samples[37850]=49754;
squeal_samples[37851]=50654;
squeal_samples[37852]=51502;
squeal_samples[37853]=52323;
squeal_samples[37854]=53101;
squeal_samples[37855]=53853;
squeal_samples[37856]=54558;
squeal_samples[37857]=52643;
squeal_samples[37858]=46784;
squeal_samples[37859]=41256;
squeal_samples[37860]=36072;
squeal_samples[37861]=31229;
squeal_samples[37862]=26691;
squeal_samples[37863]=22442;
squeal_samples[37864]=18467;
squeal_samples[37865]=14752;
squeal_samples[37866]=11276;
squeal_samples[37867]=8018;
squeal_samples[37868]=4967;
squeal_samples[37869]=4327;
squeal_samples[37870]=7199;
squeal_samples[37871]=9985;
squeal_samples[37872]=12662;
squeal_samples[37873]=15209;
squeal_samples[37874]=17653;
squeal_samples[37875]=19977;
squeal_samples[37876]=22212;
squeal_samples[37877]=24338;
squeal_samples[37878]=26373;
squeal_samples[37879]=28321;
squeal_samples[37880]=30178;
squeal_samples[37881]=31952;
squeal_samples[37882]=33651;
squeal_samples[37883]=35266;
squeal_samples[37884]=36814;
squeal_samples[37885]=38288;
squeal_samples[37886]=39701;
squeal_samples[37887]=41051;
squeal_samples[37888]=42334;
squeal_samples[37889]=43567;
squeal_samples[37890]=44730;
squeal_samples[37891]=45862;
squeal_samples[37892]=46925;
squeal_samples[37893]=47948;
squeal_samples[37894]=48926;
squeal_samples[37895]=49857;
squeal_samples[37896]=50751;
squeal_samples[37897]=51596;
squeal_samples[37898]=52413;
squeal_samples[37899]=53186;
squeal_samples[37900]=53926;
squeal_samples[37901]=54638;
squeal_samples[37902]=52711;
squeal_samples[37903]=46852;
squeal_samples[37904]=41318;
squeal_samples[37905]=36129;
squeal_samples[37906]=31282;
squeal_samples[37907]=26737;
squeal_samples[37908]=22489;
squeal_samples[37909]=18512;
squeal_samples[37910]=14789;
squeal_samples[37911]=11310;
squeal_samples[37912]=8050;
squeal_samples[37913]=5001;
squeal_samples[37914]=4353;
squeal_samples[37915]=7223;
squeal_samples[37916]=10006;
squeal_samples[37917]=12684;
squeal_samples[37918]=15227;
squeal_samples[37919]=17674;
squeal_samples[37920]=19994;
squeal_samples[37921]=22229;
squeal_samples[37922]=24353;
squeal_samples[37923]=26391;
squeal_samples[37924]=28333;
squeal_samples[37925]=30188;
squeal_samples[37926]=31964;
squeal_samples[37927]=33656;
squeal_samples[37928]=35276;
squeal_samples[37929]=36828;
squeal_samples[37930]=38297;
squeal_samples[37931]=39709;
squeal_samples[37932]=41054;
squeal_samples[37933]=42343;
squeal_samples[37934]=43570;
squeal_samples[37935]=44738;
squeal_samples[37936]=45861;
squeal_samples[37937]=46926;
squeal_samples[37938]=47955;
squeal_samples[37939]=48924;
squeal_samples[37940]=49860;
squeal_samples[37941]=50749;
squeal_samples[37942]=51598;
squeal_samples[37943]=52409;
squeal_samples[37944]=53184;
squeal_samples[37945]=53929;
squeal_samples[37946]=54636;
squeal_samples[37947]=52712;
squeal_samples[37948]=46848;
squeal_samples[37949]=41311;
squeal_samples[37950]=36127;
squeal_samples[37951]=31275;
squeal_samples[37952]=26737;
squeal_samples[37953]=22485;
squeal_samples[37954]=18505;
squeal_samples[37955]=14787;
squeal_samples[37956]=11303;
squeal_samples[37957]=8046;
squeal_samples[37958]=4989;
squeal_samples[37959]=4344;
squeal_samples[37960]=7217;
squeal_samples[37961]=10002;
squeal_samples[37962]=12673;
squeal_samples[37963]=15221;
squeal_samples[37964]=17665;
squeal_samples[37965]=19987;
squeal_samples[37966]=22221;
squeal_samples[37967]=24341;
squeal_samples[37968]=26381;
squeal_samples[37969]=28322;
squeal_samples[37970]=30183;
squeal_samples[37971]=31954;
squeal_samples[37972]=33651;
squeal_samples[37973]=35266;
squeal_samples[37974]=36816;
squeal_samples[37975]=38289;
squeal_samples[37976]=39701;
squeal_samples[37977]=41047;
squeal_samples[37978]=42330;
squeal_samples[37979]=43559;
squeal_samples[37980]=44730;
squeal_samples[37981]=45855;
squeal_samples[37982]=46921;
squeal_samples[37983]=47944;
squeal_samples[37984]=48919;
squeal_samples[37985]=49850;
squeal_samples[37986]=50739;
squeal_samples[37987]=51587;
squeal_samples[37988]=52404;
squeal_samples[37989]=53174;
squeal_samples[37990]=53918;
squeal_samples[37991]=54626;
squeal_samples[37992]=52702;
squeal_samples[37993]=46836;
squeal_samples[37994]=41304;
squeal_samples[37995]=36118;
squeal_samples[37996]=31267;
squeal_samples[37997]=26726;
squeal_samples[37998]=22474;
squeal_samples[37999]=18497;
squeal_samples[38000]=14773;
squeal_samples[38001]=11296;
squeal_samples[38002]=8032;
squeal_samples[38003]=4982;
squeal_samples[38004]=4332;
squeal_samples[38005]=7206;
squeal_samples[38006]=9993;
squeal_samples[38007]=12661;
squeal_samples[38008]=15211;
squeal_samples[38009]=17656;
squeal_samples[38010]=19975;
squeal_samples[38011]=22211;
squeal_samples[38012]=24330;
squeal_samples[38013]=26372;
squeal_samples[38014]=28310;
squeal_samples[38015]=30175;
squeal_samples[38016]=31946;
squeal_samples[38017]=33642;
squeal_samples[38018]=35256;
squeal_samples[38019]=36805;
squeal_samples[38020]=38279;
squeal_samples[38021]=39690;
squeal_samples[38022]=41036;
squeal_samples[38023]=42321;
squeal_samples[38024]=43549;
squeal_samples[38025]=44718;
squeal_samples[38026]=45844;
squeal_samples[38027]=46912;
squeal_samples[38028]=47933;
squeal_samples[38029]=48910;
squeal_samples[38030]=49837;
squeal_samples[38031]=50731;
squeal_samples[38032]=51574;
squeal_samples[38033]=52395;
squeal_samples[38034]=53163;
squeal_samples[38035]=53908;
squeal_samples[38036]=54616;
squeal_samples[38037]=52690;
squeal_samples[38038]=46828;
squeal_samples[38039]=41289;
squeal_samples[38040]=36114;
squeal_samples[38041]=31251;
squeal_samples[38042]=26719;
squeal_samples[38043]=22462;
squeal_samples[38044]=18486;
squeal_samples[38045]=14765;
squeal_samples[38046]=11282;
squeal_samples[38047]=8026;
squeal_samples[38048]=4968;
squeal_samples[38049]=4323;
squeal_samples[38050]=7196;
squeal_samples[38051]=9980;
squeal_samples[38052]=12654;
squeal_samples[38053]=15200;
squeal_samples[38054]=17642;
squeal_samples[38055]=19970;
squeal_samples[38056]=22195;
squeal_samples[38057]=24324;
squeal_samples[38058]=26360;
squeal_samples[38059]=28299;
squeal_samples[38060]=30165;
squeal_samples[38061]=31936;
squeal_samples[38062]=33631;
squeal_samples[38063]=35247;
squeal_samples[38064]=36793;
squeal_samples[38065]=38269;
squeal_samples[38066]=39681;
squeal_samples[38067]=41024;
squeal_samples[38068]=42312;
squeal_samples[38069]=43537;
squeal_samples[38070]=44710;
squeal_samples[38071]=45832;
squeal_samples[38072]=46903;
squeal_samples[38073]=47920;
squeal_samples[38074]=48902;
squeal_samples[38075]=49826;
squeal_samples[38076]=50720;
squeal_samples[38077]=51566;
squeal_samples[38078]=52381;
squeal_samples[38079]=53156;
squeal_samples[38080]=53895;
squeal_samples[38081]=54607;
squeal_samples[38082]=52680;
squeal_samples[38083]=46815;
squeal_samples[38084]=41283;
squeal_samples[38085]=36097;
squeal_samples[38086]=31248;
squeal_samples[38087]=26703;
squeal_samples[38088]=22456;
squeal_samples[38089]=18472;
squeal_samples[38090]=14756;
squeal_samples[38091]=11272;
squeal_samples[38092]=8014;
squeal_samples[38093]=4960;
squeal_samples[38094]=4312;
squeal_samples[38095]=7183;
squeal_samples[38096]=9975;
squeal_samples[38097]=12637;
squeal_samples[38098]=15195;
squeal_samples[38099]=17629;
squeal_samples[38100]=19960;
squeal_samples[38101]=22185;
squeal_samples[38102]=24314;
squeal_samples[38103]=26347;
squeal_samples[38104]=28292;
squeal_samples[38105]=30153;
squeal_samples[38106]=31926;
squeal_samples[38107]=33620;
squeal_samples[38108]=35236;
squeal_samples[38109]=36784;
squeal_samples[38110]=38258;
squeal_samples[38111]=39671;
squeal_samples[38112]=41012;
squeal_samples[38113]=42303;
squeal_samples[38114]=43526;
squeal_samples[38115]=44699;
squeal_samples[38116]=45823;
squeal_samples[38117]=46890;
squeal_samples[38118]=47913;
squeal_samples[38119]=48889;
squeal_samples[38120]=49817;
squeal_samples[38121]=50709;
squeal_samples[38122]=51555;
squeal_samples[38123]=52372;
squeal_samples[38124]=53144;
squeal_samples[38125]=53886;
squeal_samples[38126]=54596;
squeal_samples[38127]=52669;
squeal_samples[38128]=46808;
squeal_samples[38129]=41267;
squeal_samples[38130]=36092;
squeal_samples[38131]=31233;
squeal_samples[38132]=26696;
squeal_samples[38133]=22444;
squeal_samples[38134]=18463;
squeal_samples[38135]=14743;
squeal_samples[38136]=11265;
squeal_samples[38137]=8000;
squeal_samples[38138]=4954;
squeal_samples[38139]=4295;
squeal_samples[38140]=7181;
squeal_samples[38141]=9956;
squeal_samples[38142]=12634;
squeal_samples[38143]=15179;
squeal_samples[38144]=17623;
squeal_samples[38145]=19946;
squeal_samples[38146]=22178;
squeal_samples[38147]=24301;
squeal_samples[38148]=26339;
squeal_samples[38149]=28280;
squeal_samples[38150]=30143;
squeal_samples[38151]=31914;
squeal_samples[38152]=33613;
squeal_samples[38153]=35223;
squeal_samples[38154]=36775;
squeal_samples[38155]=38247;
squeal_samples[38156]=39659;
squeal_samples[38157]=41004;
squeal_samples[38158]=42291;
squeal_samples[38159]=43516;
squeal_samples[38160]=44690;
squeal_samples[38161]=45811;
squeal_samples[38162]=46880;
squeal_samples[38163]=47903;
squeal_samples[38164]=48876;
squeal_samples[38165]=49810;
squeal_samples[38166]=50697;
squeal_samples[38167]=51545;
squeal_samples[38168]=52361;
squeal_samples[38169]=53135;
squeal_samples[38170]=53872;
squeal_samples[38171]=54590;
squeal_samples[38172]=52656;
squeal_samples[38173]=46797;
squeal_samples[38174]=41260;
squeal_samples[38175]=36077;
squeal_samples[38176]=31227;
squeal_samples[38177]=26681;
squeal_samples[38178]=22438;
squeal_samples[38179]=18448;
squeal_samples[38180]=14737;
squeal_samples[38181]=11251;
squeal_samples[38182]=7992;
squeal_samples[38183]=4941;
squeal_samples[38184]=4288;
squeal_samples[38185]=7166;
squeal_samples[38186]=9950;
squeal_samples[38187]=12621;
squeal_samples[38188]=15169;
squeal_samples[38189]=17613;
squeal_samples[38190]=19936;
squeal_samples[38191]=22165;
squeal_samples[38192]=24294;
squeal_samples[38193]=26325;
squeal_samples[38194]=28273;
squeal_samples[38195]=30130;
squeal_samples[38196]=31906;
squeal_samples[38197]=33598;
squeal_samples[38198]=35218;
squeal_samples[38199]=36760;
squeal_samples[38200]=38240;
squeal_samples[38201]=39647;
squeal_samples[38202]=40993;
squeal_samples[38203]=42282;
squeal_samples[38204]=43504;
squeal_samples[38205]=44680;
squeal_samples[38206]=45801;
squeal_samples[38207]=46870;
squeal_samples[38208]=47891;
squeal_samples[38209]=48868;
squeal_samples[38210]=49795;
squeal_samples[38211]=50690;
squeal_samples[38212]=51532;
squeal_samples[38213]=52354;
squeal_samples[38214]=53118;
squeal_samples[38215]=53868;
squeal_samples[38216]=54572;
squeal_samples[38217]=53335;
squeal_samples[38218]=47582;
squeal_samples[38219]=41995;
squeal_samples[38220]=36761;
squeal_samples[38221]=31868;
squeal_samples[38222]=27280;
squeal_samples[38223]=22994;
squeal_samples[38224]=18975;
squeal_samples[38225]=15222;
squeal_samples[38226]=11709;
squeal_samples[38227]=8417;
squeal_samples[38228]=5340;
squeal_samples[38229]=4087;
squeal_samples[38230]=6831;
squeal_samples[38231]=9637;
squeal_samples[38232]=12315;
squeal_samples[38233]=14880;
squeal_samples[38234]=17331;
squeal_samples[38235]=19670;
squeal_samples[38236]=21907;
squeal_samples[38237]=24051;
squeal_samples[38238]=26094;
squeal_samples[38239]=28047;
squeal_samples[38240]=29916;
squeal_samples[38241]=31694;
squeal_samples[38242]=33399;
squeal_samples[38243]=35026;
squeal_samples[38244]=36584;
squeal_samples[38245]=38063;
squeal_samples[38246]=39482;
squeal_samples[38247]=40837;
squeal_samples[38248]=42127;
squeal_samples[38249]=43362;
squeal_samples[38250]=44540;
squeal_samples[38251]=45668;
squeal_samples[38252]=46741;
squeal_samples[38253]=47765;
squeal_samples[38254]=48751;
squeal_samples[38255]=49679;
squeal_samples[38256]=50583;
squeal_samples[38257]=51430;
squeal_samples[38258]=52248;
squeal_samples[38259]=53026;
squeal_samples[38260]=53770;
squeal_samples[38261]=54489;
squeal_samples[38262]=53832;
squeal_samples[38263]=48309;
squeal_samples[38264]=42664;
squeal_samples[38265]=37398;
squeal_samples[38266]=32453;
squeal_samples[38267]=27841;
squeal_samples[38268]=23505;
squeal_samples[38269]=19462;
squeal_samples[38270]=15670;
squeal_samples[38271]=12130;
squeal_samples[38272]=8814;
squeal_samples[38273]=5705;
squeal_samples[38274]=3934;
squeal_samples[38275]=6461;
squeal_samples[38276]=9285;
squeal_samples[38277]=11980;
squeal_samples[38278]=14557;
squeal_samples[38279]=17026;
squeal_samples[38280]=19373;
squeal_samples[38281]=21630;
squeal_samples[38282]=23776;
squeal_samples[38283]=25836;
squeal_samples[38284]=27796;
squeal_samples[38285]=29680;
squeal_samples[38286]=31471;
squeal_samples[38287]=33182;
squeal_samples[38288]=34822;
squeal_samples[38289]=36381;
squeal_samples[38290]=37877;
squeal_samples[38291]=39301;
squeal_samples[38292]=40658;
squeal_samples[38293]=41962;
squeal_samples[38294]=43201;
squeal_samples[38295]=44389;
squeal_samples[38296]=45517;
squeal_samples[38297]=46602;
squeal_samples[38298]=47630;
squeal_samples[38299]=48619;
squeal_samples[38300]=49559;
squeal_samples[38301]=50459;
squeal_samples[38302]=51320;
squeal_samples[38303]=52138;
squeal_samples[38304]=52923;
squeal_samples[38305]=53673;
squeal_samples[38306]=54390;
squeal_samples[38307]=54220;
squeal_samples[38308]=49025;
squeal_samples[38309]=43339;
squeal_samples[38310]=38028;
squeal_samples[38311]=33040;
squeal_samples[38312]=28390;
squeal_samples[38313]=24021;
squeal_samples[38314]=19946;
squeal_samples[38315]=16122;
squeal_samples[38316]=12554;
squeal_samples[38317]=9203;
squeal_samples[38318]=6079;
squeal_samples[38319]=3864;
squeal_samples[38320]=6098;
squeal_samples[38321]=8922;
squeal_samples[38322]=11639;
squeal_samples[38323]=14235;
squeal_samples[38324]=16706;
squeal_samples[38325]=19079;
squeal_samples[38326]=21341;
squeal_samples[38327]=23504;
squeal_samples[38328]=25579;
squeal_samples[38329]=27546;
squeal_samples[38330]=29439;
squeal_samples[38331]=31242;
squeal_samples[38332]=32961;
squeal_samples[38333]=34614;
squeal_samples[38334]=36179;
squeal_samples[38335]=37683;
squeal_samples[38336]=39112;
squeal_samples[38337]=40484;
squeal_samples[38338]=41794;
squeal_samples[38339]=43040;
squeal_samples[38340]=44230;
squeal_samples[38341]=45368;
squeal_samples[38342]=46459;
squeal_samples[38343]=47497;
squeal_samples[38344]=48488;
squeal_samples[38345]=49435;
squeal_samples[38346]=50340;
squeal_samples[38347]=51206;
squeal_samples[38348]=52024;
squeal_samples[38349]=52816;
squeal_samples[38350]=53569;
squeal_samples[38351]=54292;
squeal_samples[38352]=54499;
squeal_samples[38353]=49749;
squeal_samples[38354]=44027;
squeal_samples[38355]=38654;
squeal_samples[38356]=33647;
squeal_samples[38357]=28937;
squeal_samples[38358]=24543;
squeal_samples[38359]=20424;
squeal_samples[38360]=16585;
squeal_samples[38361]=12971;
squeal_samples[38362]=9608;
squeal_samples[38363]=6441;
squeal_samples[38364]=3905;
squeal_samples[38365]=5716;
squeal_samples[38366]=8570;
squeal_samples[38367]=11293;
squeal_samples[38368]=13904;
squeal_samples[38369]=16396;
squeal_samples[38370]=18770;
squeal_samples[38371]=21058;
squeal_samples[38372]=23227;
squeal_samples[38373]=25311;
squeal_samples[38374]=27295;
squeal_samples[38375]=29193;
squeal_samples[38376]=31008;
squeal_samples[38377]=32745;
squeal_samples[38378]=34395;
squeal_samples[38379]=35981;
squeal_samples[38380]=37482;
squeal_samples[38381]=38930;
squeal_samples[38382]=40307;
squeal_samples[38383]=41619;
squeal_samples[38384]=42879;
squeal_samples[38385]=44077;
squeal_samples[38386]=45222;
squeal_samples[38387]=46315;
squeal_samples[38388]=47359;
squeal_samples[38389]=48356;
squeal_samples[38390]=49308;
squeal_samples[38391]=50217;
squeal_samples[38392]=51086;
squeal_samples[38393]=51917;
squeal_samples[38394]=52711;
squeal_samples[38395]=53470;
squeal_samples[38396]=54191;
squeal_samples[38397]=54673;
squeal_samples[38398]=50486;
squeal_samples[38399]=44707;
squeal_samples[38400]=39301;
squeal_samples[38401]=34240;
squeal_samples[38402]=29500;
squeal_samples[38403]=25068;
squeal_samples[38404]=20916;
squeal_samples[38405]=17038;
squeal_samples[38406]=13399;
squeal_samples[38407]=10001;
squeal_samples[38408]=6815;
squeal_samples[38409]=4022;
squeal_samples[38410]=5344;
squeal_samples[38411]=8209;
squeal_samples[38412]=10955;
squeal_samples[38413]=13569;
squeal_samples[38414]=16084;
squeal_samples[38415]=18468;
squeal_samples[38416]=20761;
squeal_samples[38417]=22955;
squeal_samples[38418]=25042;
squeal_samples[38419]=27047;
squeal_samples[38420]=28950;
squeal_samples[38421]=30782;
squeal_samples[38422]=32518;
squeal_samples[38423]=34186;
squeal_samples[38424]=35767;
squeal_samples[38425]=37294;
squeal_samples[38426]=38737;
squeal_samples[38427]=40131;
squeal_samples[38428]=41444;
squeal_samples[38429]=42712;
squeal_samples[38430]=43915;
squeal_samples[38431]=45071;
squeal_samples[38432]=46168;
squeal_samples[38433]=47220;
squeal_samples[38434]=48224;
squeal_samples[38435]=49181;
squeal_samples[38436]=50096;
squeal_samples[38437]=50973;
squeal_samples[38438]=51804;
squeal_samples[38439]=52602;
squeal_samples[38440]=53367;
squeal_samples[38441]=54089;
squeal_samples[38442]=54736;
squeal_samples[38443]=51223;
squeal_samples[38444]=45401;
squeal_samples[38445]=39949;
squeal_samples[38446]=34843;
squeal_samples[38447]=30065;
squeal_samples[38448]=25595;
squeal_samples[38449]=21412;
squeal_samples[38450]=17498;
squeal_samples[38451]=13836;
squeal_samples[38452]=10402;
squeal_samples[38453]=7192;
squeal_samples[38454]=4233;
squeal_samples[38455]=4971;
squeal_samples[38456]=7848;
squeal_samples[38457]=10610;
squeal_samples[38458]=13239;
squeal_samples[38459]=15762;
squeal_samples[38460]=18172;
squeal_samples[38461]=20472;
squeal_samples[38462]=22674;
squeal_samples[38463]=24777;
squeal_samples[38464]=26787;
squeal_samples[38465]=28707;
squeal_samples[38466]=30542;
squeal_samples[38467]=32292;
squeal_samples[38468]=33974;
squeal_samples[38469]=35563;
squeal_samples[38470]=37098;
squeal_samples[38471]=38554;
squeal_samples[38472]=39945;
squeal_samples[38473]=41278;
squeal_samples[38474]=42550;
squeal_samples[38475]=43757;
squeal_samples[38476]=44921;
squeal_samples[38477]=46026;
squeal_samples[38478]=47079;
squeal_samples[38479]=48090;
squeal_samples[38480]=49055;
squeal_samples[38481]=49973;
squeal_samples[38482]=50854;
squeal_samples[38483]=51689;
squeal_samples[38484]=52495;
squeal_samples[38485]=53263;
squeal_samples[38486]=53992;
squeal_samples[38487]=54693;
squeal_samples[38488]=51967;
squeal_samples[38489]=46097;
squeal_samples[38490]=40602;
squeal_samples[38491]=35452;
squeal_samples[38492]=30634;
squeal_samples[38493]=26130;
squeal_samples[38494]=21909;
squeal_samples[38495]=17963;
squeal_samples[38496]=14264;
squeal_samples[38497]=10810;
squeal_samples[38498]=7572;
squeal_samples[38499]=4546;
squeal_samples[38500]=4587;
squeal_samples[38501]=7489;
squeal_samples[38502]=10259;
squeal_samples[38503]=12909;
squeal_samples[38504]=15448;
squeal_samples[38505]=17867;
squeal_samples[38506]=20182;
squeal_samples[38507]=22395;
squeal_samples[38508]=24509;
squeal_samples[38509]=26529;
squeal_samples[38510]=28466;
squeal_samples[38511]=30306;
squeal_samples[38512]=32075;
squeal_samples[38513]=33752;
squeal_samples[38514]=35362;
squeal_samples[38515]=36894;
squeal_samples[38516]=38367;
squeal_samples[38517]=39765;
squeal_samples[38518]=41106;
squeal_samples[38519]=42382;
squeal_samples[38520]=43600;
squeal_samples[38521]=44770;
squeal_samples[38522]=45880;
squeal_samples[38523]=46938;
squeal_samples[38524]=47956;
squeal_samples[38525]=48923;
squeal_samples[38526]=49852;
squeal_samples[38527]=50731;
squeal_samples[38528]=51580;
squeal_samples[38529]=52382;
squeal_samples[38530]=53157;
squeal_samples[38531]=53894;
squeal_samples[38532]=54600;
squeal_samples[38533]=52670;
squeal_samples[38534]=46796;
squeal_samples[38535]=41262;
squeal_samples[38536]=36063;
squeal_samples[38537]=31215;
squeal_samples[38538]=26664;
squeal_samples[38539]=22411;
squeal_samples[38540]=18424;
squeal_samples[38541]=14705;
squeal_samples[38542]=11219;
squeal_samples[38543]=7952;
squeal_samples[38544]=4904;
squeal_samples[38545]=4252;
squeal_samples[38546]=7119;
squeal_samples[38547]=9907;
squeal_samples[38548]=12573;
squeal_samples[38549]=15121;
squeal_samples[38550]=17560;
squeal_samples[38551]=19882;
squeal_samples[38552]=22117;
squeal_samples[38553]=24237;
squeal_samples[38554]=26277;
squeal_samples[38555]=28210;
squeal_samples[38556]=30073;
squeal_samples[38557]=31844;
squeal_samples[38558]=33537;
squeal_samples[38559]=35156;
squeal_samples[38560]=36699;
squeal_samples[38561]=38177;
squeal_samples[38562]=39583;
squeal_samples[38563]=40926;
squeal_samples[38564]=42213;
squeal_samples[38565]=43441;
squeal_samples[38566]=44608;
squeal_samples[38567]=45739;
squeal_samples[38568]=46794;
squeal_samples[38569]=47822;
squeal_samples[38570]=48793;
squeal_samples[38571]=49727;
squeal_samples[38572]=50612;
squeal_samples[38573]=51465;
squeal_samples[38574]=52276;
squeal_samples[38575]=53052;
squeal_samples[38576]=53790;
squeal_samples[38577]=54503;
squeal_samples[38578]=53841;
squeal_samples[38579]=48311;
squeal_samples[38580]=42670;
squeal_samples[38581]=37394;
squeal_samples[38582]=32447;
squeal_samples[38583]=27827;
squeal_samples[38584]=23487;
squeal_samples[38585]=19444;
squeal_samples[38586]=15647;
squeal_samples[38587]=12106;
squeal_samples[38588]=8784;
squeal_samples[38589]=5676;
squeal_samples[38590]=3900;
squeal_samples[38591]=6427;
squeal_samples[38592]=9245;
squeal_samples[38593]=11938;
squeal_samples[38594]=14520;
squeal_samples[38595]=16977;
squeal_samples[38596]=19333;
squeal_samples[38597]=21579;
squeal_samples[38598]=23735;
squeal_samples[38599]=25787;
squeal_samples[38600]=27755;
squeal_samples[38601]=29626;
squeal_samples[38602]=31421;
squeal_samples[38603]=33132;
squeal_samples[38604]=34769;
squeal_samples[38605]=36329;
squeal_samples[38606]=37815;
squeal_samples[38607]=39251;
squeal_samples[38608]=40597;
squeal_samples[38609]=41909;
squeal_samples[38610]=43144;
squeal_samples[38611]=44331;
squeal_samples[38612]=45457;
squeal_samples[38613]=46539;
squeal_samples[38614]=47575;
squeal_samples[38615]=48557;
squeal_samples[38616]=49498;
squeal_samples[38617]=50396;
squeal_samples[38618]=51258;
squeal_samples[38619]=52076;
squeal_samples[38620]=52862;
squeal_samples[38621]=53606;
squeal_samples[38622]=54327;
squeal_samples[38623]=54528;
squeal_samples[38624]=49776;
squeal_samples[38625]=44042;
squeal_samples[38626]=38672;
squeal_samples[38627]=33653;
squeal_samples[38628]=28947;
squeal_samples[38629]=24545;
squeal_samples[38630]=20423;
squeal_samples[38631]=16574;
squeal_samples[38632]=12962;
squeal_samples[38633]=9585;
squeal_samples[38634]=6426;
squeal_samples[38635]=3879;
squeal_samples[38636]=5699;
squeal_samples[38637]=8544;
squeal_samples[38638]=11271;
squeal_samples[38639]=13878;
squeal_samples[38640]=16366;
squeal_samples[38641]=18745;
squeal_samples[38642]=21017;
squeal_samples[38643]=23197;
squeal_samples[38644]=25273;
squeal_samples[38645]=27260;
squeal_samples[38646]=29161;
squeal_samples[38647]=30970;
squeal_samples[38648]=32705;
squeal_samples[38649]=34357;
squeal_samples[38650]=35937;
squeal_samples[38651]=37446;
squeal_samples[38652]=38886;
squeal_samples[38653]=40264;
squeal_samples[38654]=41571;
squeal_samples[38655]=42835;
squeal_samples[38656]=44031;
squeal_samples[38657]=45170;
squeal_samples[38658]=46269;
squeal_samples[38659]=47309;
squeal_samples[38660]=48308;
squeal_samples[38661]=49259;
squeal_samples[38662]=50165;
squeal_samples[38663]=51033;
squeal_samples[38664]=51868;
squeal_samples[38665]=52658;
squeal_samples[38666]=53418;
squeal_samples[38667]=54141;
squeal_samples[38668]=54776;
squeal_samples[38669]=51264;
squeal_samples[38670]=45431;
squeal_samples[38671]=39972;
squeal_samples[38672]=34863;
squeal_samples[38673]=30081;
squeal_samples[38674]=25613;
squeal_samples[38675]=21415;
squeal_samples[38676]=17505;
squeal_samples[38677]=13830;
squeal_samples[38678]=10400;
squeal_samples[38679]=7188;
squeal_samples[38680]=4227;
squeal_samples[38681]=4954;
squeal_samples[38682]=7839;
squeal_samples[38683]=10592;
squeal_samples[38684]=13227;
squeal_samples[38685]=15748;
squeal_samples[38686]=18153;
squeal_samples[38687]=20448;
squeal_samples[38688]=22654;
squeal_samples[38689]=24753;
squeal_samples[38690]=26762;
squeal_samples[38691]=28683;
squeal_samples[38692]=30517;
squeal_samples[38693]=32268;
squeal_samples[38694]=33943;
squeal_samples[38695]=35533;
squeal_samples[38696]=37069;
squeal_samples[38697]=38518;
squeal_samples[38698]=39914;
squeal_samples[38699]=41245;
squeal_samples[38700]=42511;
squeal_samples[38701]=43726;
squeal_samples[38702]=44882;
squeal_samples[38703]=45987;
squeal_samples[38704]=47043;
squeal_samples[38705]=48055;
squeal_samples[38706]=49013;
squeal_samples[38707]=49934;
squeal_samples[38708]=50811;
squeal_samples[38709]=51650;
squeal_samples[38710]=52452;
squeal_samples[38711]=53223;
squeal_samples[38712]=53950;
squeal_samples[38713]=54651;
squeal_samples[38714]=52715;
squeal_samples[38715]=46838;
squeal_samples[38716]=41294;
squeal_samples[38717]=36101;
squeal_samples[38718]=31240;
squeal_samples[38719]=26691;
squeal_samples[38720]=22428;
squeal_samples[38721]=18443;
squeal_samples[38722]=14718;
squeal_samples[38723]=11225;
squeal_samples[38724]=7962;
squeal_samples[38725]=4899;
squeal_samples[38726]=4250;
squeal_samples[38727]=7115;
squeal_samples[38728]=9903;
squeal_samples[38729]=12566;
squeal_samples[38730]=15117;
squeal_samples[38731]=17551;
squeal_samples[38732]=19874;
squeal_samples[38733]=22100;
squeal_samples[38734]=24229;
squeal_samples[38735]=26256;
squeal_samples[38736]=28201;
squeal_samples[38737]=30057;
squeal_samples[38738]=31823;
squeal_samples[38739]=33520;
squeal_samples[38740]=35135;
squeal_samples[38741]=36679;
squeal_samples[38742]=38156;
squeal_samples[38743]=39557;
squeal_samples[38744]=40911;
squeal_samples[38745]=42188;
squeal_samples[38746]=43413;
squeal_samples[38747]=44588;
squeal_samples[38748]=45703;
squeal_samples[38749]=46773;
squeal_samples[38750]=47796;
squeal_samples[38751]=48763;
squeal_samples[38752]=49700;
squeal_samples[38753]=50585;
squeal_samples[38754]=51431;
squeal_samples[38755]=52250;
squeal_samples[38756]=53018;
squeal_samples[38757]=53762;
squeal_samples[38758]=54471;
squeal_samples[38759]=53812;
squeal_samples[38760]=48276;
squeal_samples[38761]=42632;
squeal_samples[38762]=37360;
squeal_samples[38763]=32410;
squeal_samples[38764]=27792;
squeal_samples[38765]=23453;
squeal_samples[38766]=19404;
squeal_samples[38767]=15616;
squeal_samples[38768]=12066;
squeal_samples[38769]=8746;
squeal_samples[38770]=5639;
squeal_samples[38771]=3864;
squeal_samples[38772]=6392;
squeal_samples[38773]=9209;
squeal_samples[38774]=11903;
squeal_samples[38775]=14477;
squeal_samples[38776]=16943;
squeal_samples[38777]=19296;
squeal_samples[38778]=21539;
squeal_samples[38779]=23699;
squeal_samples[38780]=25746;
squeal_samples[38781]=27713;
squeal_samples[38782]=29591;
squeal_samples[38783]=31380;
squeal_samples[38784]=33096;
squeal_samples[38785]=34729;
squeal_samples[38786]=36290;
squeal_samples[38787]=37785;
squeal_samples[38788]=39204;
squeal_samples[38789]=40566;
squeal_samples[38790]=41864;
squeal_samples[38791]=43104;
squeal_samples[38792]=44290;
squeal_samples[38793]=45423;
squeal_samples[38794]=46501;
squeal_samples[38795]=47535;
squeal_samples[38796]=48515;
squeal_samples[38797]=49462;
squeal_samples[38798]=50356;
squeal_samples[38799]=51217;
squeal_samples[38800]=52034;
squeal_samples[38801]=52822;
squeal_samples[38802]=53569;
squeal_samples[38803]=54286;
squeal_samples[38804]=54488;
squeal_samples[38805]=49734;
squeal_samples[38806]=44002;
squeal_samples[38807]=38631;
squeal_samples[38808]=33610;
squeal_samples[38809]=28908;
squeal_samples[38810]=24502;
squeal_samples[38811]=20384;
squeal_samples[38812]=16531;
squeal_samples[38813]=12923;
squeal_samples[38814]=9542;
squeal_samples[38815]=6386;
squeal_samples[38816]=3837;
squeal_samples[38817]=5657;
squeal_samples[38818]=8511;
squeal_samples[38819]=11227;
squeal_samples[38820]=13840;
squeal_samples[38821]=16323;
squeal_samples[38822]=18703;
squeal_samples[38823]=20984;
squeal_samples[38824]=23153;
squeal_samples[38825]=25233;
squeal_samples[38826]=27221;
squeal_samples[38827]=29116;
squeal_samples[38828]=30933;
squeal_samples[38829]=32662;
squeal_samples[38830]=34316;
squeal_samples[38831]=35896;
squeal_samples[38832]=37405;
squeal_samples[38833]=38845;
squeal_samples[38834]=40222;
squeal_samples[38835]=41532;
squeal_samples[38836]=42792;
squeal_samples[38837]=43990;
squeal_samples[38838]=45132;
squeal_samples[38839]=46223;
squeal_samples[38840]=47272;
squeal_samples[38841]=48265;
squeal_samples[38842]=49219;
squeal_samples[38843]=50122;
squeal_samples[38844]=50995;
squeal_samples[38845]=51823;
squeal_samples[38846]=52621;
squeal_samples[38847]=53374;
squeal_samples[38848]=54101;
squeal_samples[38849]=54736;
squeal_samples[38850]=51220;
squeal_samples[38851]=45392;
squeal_samples[38852]=39930;
squeal_samples[38853]=34824;
squeal_samples[38854]=30039;
squeal_samples[38855]=25572;
squeal_samples[38856]=21372;
squeal_samples[38857]=17466;
squeal_samples[38858]=13788;
squeal_samples[38859]=10360;
squeal_samples[38860]=7148;
squeal_samples[38861]=4183;
squeal_samples[38862]=4915;
squeal_samples[38863]=7797;
squeal_samples[38864]=10550;
squeal_samples[38865]=13188;
squeal_samples[38866]=15706;
squeal_samples[38867]=18111;
squeal_samples[38868]=20409;
squeal_samples[38869]=22610;
squeal_samples[38870]=24715;
squeal_samples[38871]=26717;
squeal_samples[38872]=28646;
squeal_samples[38873]=30472;
squeal_samples[38874]=32231;
squeal_samples[38875]=33898;
squeal_samples[38876]=35495;
squeal_samples[38877]=37026;
squeal_samples[38878]=38476;
squeal_samples[38879]=39877;
squeal_samples[38880]=41199;
squeal_samples[38881]=42475;
squeal_samples[38882]=43679;
squeal_samples[38883]=44845;
squeal_samples[38884]=45944;
squeal_samples[38885]=47003;
squeal_samples[38886]=48013;
squeal_samples[38887]=48972;
squeal_samples[38888]=49892;
squeal_samples[38889]=50771;
squeal_samples[38890]=51607;
squeal_samples[38891]=52414;
squeal_samples[38892]=53177;
squeal_samples[38893]=53913;
squeal_samples[38894]=54605;
squeal_samples[38895]=53362;
squeal_samples[38896]=47593;
squeal_samples[38897]=41999;
squeal_samples[38898]=36753;
squeal_samples[38899]=31851;
squeal_samples[38900]=27258;
squeal_samples[38901]=22957;
squeal_samples[38902]=18934;
squeal_samples[38903]=15176;
squeal_samples[38904]=11651;
squeal_samples[38905]=8355;
squeal_samples[38906]=5273;
squeal_samples[38907]=4011;
squeal_samples[38908]=6753;
squeal_samples[38909]=9553;
squeal_samples[38910]=12230;
squeal_samples[38911]=14796;
squeal_samples[38912]=17242;
squeal_samples[38913]=19579;
squeal_samples[38914]=21813;
squeal_samples[38915]=23955;
squeal_samples[38916]=25992;
squeal_samples[38917]=27949;
squeal_samples[38918]=29809;
squeal_samples[38919]=31588;
squeal_samples[38920]=33293;
squeal_samples[38921]=34914;
squeal_samples[38922]=36467;
squeal_samples[38923]=37948;
squeal_samples[38924]=39364;
squeal_samples[38925]=40714;
squeal_samples[38926]=42007;
squeal_samples[38927]=43235;
squeal_samples[38928]=44418;
squeal_samples[38929]=45542;
squeal_samples[38930]=46613;
squeal_samples[38931]=47639;
squeal_samples[38932]=48621;
squeal_samples[38933]=49553;
squeal_samples[38934]=50449;
squeal_samples[38935]=51295;
squeal_samples[38936]=52116;
squeal_samples[38937]=52891;
squeal_samples[38938]=53638;
squeal_samples[38939]=54346;
squeal_samples[38940]=54549;
squeal_samples[38941]=49791;
squeal_samples[38942]=44052;
squeal_samples[38943]=38676;
squeal_samples[38944]=33651;
squeal_samples[38945]=28938;
squeal_samples[38946]=24537;
squeal_samples[38947]=20401;
squeal_samples[38948]=16561;
squeal_samples[38949]=12935;
squeal_samples[38950]=9564;
squeal_samples[38951]=6396;
squeal_samples[38952]=3852;
squeal_samples[38953]=5663;
squeal_samples[38954]=8512;
squeal_samples[38955]=11236;
squeal_samples[38956]=13838;
squeal_samples[38957]=16335;
squeal_samples[38958]=18702;
squeal_samples[38959]=20980;
squeal_samples[38960]=23156;
squeal_samples[38961]=25229;
squeal_samples[38962]=27215;
squeal_samples[38963]=29116;
squeal_samples[38964]=30921;
squeal_samples[38965]=32653;
squeal_samples[38966]=34309;
squeal_samples[38967]=35884;
squeal_samples[38968]=37397;
squeal_samples[38969]=38832;
squeal_samples[38970]=40210;
squeal_samples[38971]=41525;
squeal_samples[38972]=42776;
squeal_samples[38973]=43971;
squeal_samples[38974]=45117;
squeal_samples[38975]=46203;
squeal_samples[38976]=47257;
squeal_samples[38977]=48245;
squeal_samples[38978]=49199;
squeal_samples[38979]=50108;
squeal_samples[38980]=50973;
squeal_samples[38981]=51805;
squeal_samples[38982]=52598;
squeal_samples[38983]=53357;
squeal_samples[38984]=54072;
squeal_samples[38985]=54772;
squeal_samples[38986]=52030;
squeal_samples[38987]=46149;
squeal_samples[38988]=40639;
squeal_samples[38989]=35485;
squeal_samples[38990]=30658;
squeal_samples[38991]=26140;
squeal_samples[38992]=21916;
squeal_samples[38993]=17963;
squeal_samples[38994]=14260;
squeal_samples[38995]=10793;
squeal_samples[38996]=7553;
squeal_samples[38997]=4517;
squeal_samples[38998]=4558;
squeal_samples[38999]=7449;
squeal_samples[39000]=10218;
squeal_samples[39001]=12866;
squeal_samples[39002]=15400;
squeal_samples[39003]=17819;
squeal_samples[39004]=20127;
squeal_samples[39005]=22344;
squeal_samples[39006]=24452;
squeal_samples[39007]=26474;
squeal_samples[39008]=28399;
squeal_samples[39009]=30243;
squeal_samples[39010]=32004;
squeal_samples[39011]=33683;
squeal_samples[39012]=35291;
squeal_samples[39013]=36825;
squeal_samples[39014]=38292;
squeal_samples[39015]=39689;
squeal_samples[39016]=41027;
squeal_samples[39017]=42298;
squeal_samples[39018]=43522;
squeal_samples[39019]=44682;
squeal_samples[39020]=45794;
squeal_samples[39021]=46860;
squeal_samples[39022]=47865;
squeal_samples[39023]=48841;
squeal_samples[39024]=49762;
squeal_samples[39025]=50643;
squeal_samples[39026]=51490;
squeal_samples[39027]=52294;
squeal_samples[39028]=53061;
squeal_samples[39029]=53799;
squeal_samples[39030]=54500;
squeal_samples[39031]=53839;
squeal_samples[39032]=48299;
squeal_samples[39033]=42654;
squeal_samples[39034]=37372;
squeal_samples[39035]=32422;
squeal_samples[39036]=27792;
squeal_samples[39037]=23459;
squeal_samples[39038]=19396;
squeal_samples[39039]=15608;
squeal_samples[39040]=12054;
squeal_samples[39041]=8733;
squeal_samples[39042]=5621;
squeal_samples[39043]=3840;
squeal_samples[39044]=6368;
squeal_samples[39045]=9186;
squeal_samples[39046]=11879;
squeal_samples[39047]=14454;
squeal_samples[39048]=16915;
squeal_samples[39049]=19262;
squeal_samples[39050]=21516;
squeal_samples[39051]=23660;
squeal_samples[39052]=25713;
squeal_samples[39053]=27680;
squeal_samples[39054]=29553;
squeal_samples[39055]=31348;
squeal_samples[39056]=33056;
squeal_samples[39057]=34687;
squeal_samples[39058]=36253;
squeal_samples[39059]=37737;
squeal_samples[39060]=39166;
squeal_samples[39061]=40520;
squeal_samples[39062]=41819;
squeal_samples[39063]=43059;
squeal_samples[39064]=44244;
squeal_samples[39065]=45373;
squeal_samples[39066]=46450;
squeal_samples[39067]=47484;
squeal_samples[39068]=48471;
squeal_samples[39069]=49409;
squeal_samples[39070]=50308;
squeal_samples[39071]=51162;
squeal_samples[39072]=51988;
squeal_samples[39073]=52766;
squeal_samples[39074]=53517;
squeal_samples[39075]=54232;
squeal_samples[39076]=54703;
squeal_samples[39077]=50505;
squeal_samples[39078]=44721;
squeal_samples[39079]=39299;
squeal_samples[39080]=34226;
squeal_samples[39081]=29483;
squeal_samples[39082]=25036;
squeal_samples[39083]=20883;
squeal_samples[39084]=16990;
squeal_samples[39085]=13350;
squeal_samples[39086]=9943;
squeal_samples[39087]=6754;
squeal_samples[39088]=3948;
squeal_samples[39089]=5271;
squeal_samples[39090]=8131;
squeal_samples[39091]=10870;
squeal_samples[39092]=13487;
squeal_samples[39093]=15994;
squeal_samples[39094]=18378;
squeal_samples[39095]=20674;
squeal_samples[39096]=22857;
squeal_samples[39097]=24950;
squeal_samples[39098]=26941;
squeal_samples[39099]=28850;
squeal_samples[39100]=30676;
squeal_samples[39101]=32408;
squeal_samples[39102]=34079;
squeal_samples[39103]=35658;
squeal_samples[39104]=37182;
squeal_samples[39105]=38626;
squeal_samples[39106]=40014;
squeal_samples[39107]=41329;
squeal_samples[39108]=42590;
squeal_samples[39109]=43792;
squeal_samples[39110]=44945;
squeal_samples[39111]=46045;
squeal_samples[39112]=47093;
squeal_samples[39113]=48098;
squeal_samples[39114]=49051;
squeal_samples[39115]=49965;
squeal_samples[39116]=50840;
squeal_samples[39117]=51670;
squeal_samples[39118]=52470;
squeal_samples[39119]=53233;
squeal_samples[39120]=53954;
squeal_samples[39121]=54660;
squeal_samples[39122]=52710;
squeal_samples[39123]=46838;
squeal_samples[39124]=41278;
squeal_samples[39125]=36083;
squeal_samples[39126]=31211;
squeal_samples[39127]=26659;
squeal_samples[39128]=22396;
squeal_samples[39129]=18403;
squeal_samples[39130]=14682;
squeal_samples[39131]=11181;
squeal_samples[39132]=7911;
squeal_samples[39133]=4855;
squeal_samples[39134]=4196;
squeal_samples[39135]=7070;
squeal_samples[39136]=9846;
squeal_samples[39137]=12512;
squeal_samples[39138]=15059;
squeal_samples[39139]=17489;
squeal_samples[39140]=19818;
squeal_samples[39141]=22036;
squeal_samples[39142]=24167;
squeal_samples[39143]=26188;
squeal_samples[39144]=28138;
squeal_samples[39145]=29985;
squeal_samples[39146]=31760;
squeal_samples[39147]=33448;
squeal_samples[39148]=35064;
squeal_samples[39149]=36604;
squeal_samples[39150]=38084;
squeal_samples[39151]=39483;
squeal_samples[39152]=40835;
squeal_samples[39153]=42115;
squeal_samples[39154]=43340;
squeal_samples[39155]=44510;
squeal_samples[39156]=45628;
squeal_samples[39157]=46698;
squeal_samples[39158]=47711;
squeal_samples[39159]=48691;
squeal_samples[39160]=49616;
squeal_samples[39161]=50505;
squeal_samples[39162]=51355;
squeal_samples[39163]=52166;
squeal_samples[39164]=52939;
squeal_samples[39165]=53678;
squeal_samples[39166]=54386;
squeal_samples[39167]=54201;
squeal_samples[39168]=49005;
squeal_samples[39169]=43306;
squeal_samples[39170]=37982;
squeal_samples[39171]=32990;
squeal_samples[39172]=28320;
squeal_samples[39173]=23955;
squeal_samples[39174]=19859;
squeal_samples[39175]=16040;
squeal_samples[39176]=12451;
squeal_samples[39177]=9106;
squeal_samples[39178]=5964;
squeal_samples[39179]=3762;
squeal_samples[39180]=5977;
squeal_samples[39181]=8808;
squeal_samples[39182]=11518;
squeal_samples[39183]=14107;
squeal_samples[39184]=16587;
squeal_samples[39185]=18938;
squeal_samples[39186]=21208;
squeal_samples[39187]=23364;
squeal_samples[39188]=25433;
squeal_samples[39189]=27410;
squeal_samples[39190]=29290;
squeal_samples[39191]=31095;
squeal_samples[39192]=32812;
squeal_samples[39193]=34458;
squeal_samples[39194]=36026;
squeal_samples[39195]=37527;
squeal_samples[39196]=38956;
squeal_samples[39197]=40322;
squeal_samples[39198]=41630;
squeal_samples[39199]=42879;
squeal_samples[39200]=44064;
squeal_samples[39201]=45207;
squeal_samples[39202]=46290;
squeal_samples[39203]=47329;
squeal_samples[39204]=48319;
squeal_samples[39205]=49268;
squeal_samples[39206]=50164;
squeal_samples[39207]=51033;
squeal_samples[39208]=51856;
squeal_samples[39209]=52640;
squeal_samples[39210]=53397;
squeal_samples[39211]=54110;
squeal_samples[39212]=54753;
squeal_samples[39213]=51225;
squeal_samples[39214]=45391;
squeal_samples[39215]=39924;
squeal_samples[39216]=34817;
squeal_samples[39217]=30024;
squeal_samples[39218]=25548;
squeal_samples[39219]=21353;
squeal_samples[39220]=17435;
squeal_samples[39221]=13763;
squeal_samples[39222]=10325;
squeal_samples[39223]=7110;
squeal_samples[39224]=4146;
squeal_samples[39225]=4870;
squeal_samples[39226]=7754;
squeal_samples[39227]=10500;
squeal_samples[39228]=13140;
squeal_samples[39229]=15653;
squeal_samples[39230]=18061;
squeal_samples[39231]=20356;
squeal_samples[39232]=22559;
squeal_samples[39233]=24656;
squeal_samples[39234]=26666;
squeal_samples[39235]=28588;
squeal_samples[39236]=30414;
squeal_samples[39237]=32171;
squeal_samples[39238]=33836;
squeal_samples[39239]=35437;
squeal_samples[39240]=36958;
squeal_samples[39241]=38419;
squeal_samples[39242]=39808;
squeal_samples[39243]=41136;
squeal_samples[39244]=42407;
squeal_samples[39245]=43616;
squeal_samples[39246]=44773;
squeal_samples[39247]=45877;
squeal_samples[39248]=46934;
squeal_samples[39249]=47940;
squeal_samples[39250]=48903;
squeal_samples[39251]=49825;
squeal_samples[39252]=50700;
squeal_samples[39253]=51536;
squeal_samples[39254]=52341;
squeal_samples[39255]=53104;
squeal_samples[39256]=53836;
squeal_samples[39257]=54540;
squeal_samples[39258]=53866;
squeal_samples[39259]=48324;
squeal_samples[39260]=42676;
squeal_samples[39261]=37383;
squeal_samples[39262]=32432;
squeal_samples[39263]=27802;
squeal_samples[39264]=23458;
squeal_samples[39265]=19404;
squeal_samples[39266]=15602;
squeal_samples[39267]=12049;
squeal_samples[39268]=8723;
squeal_samples[39269]=5610;
squeal_samples[39270]=3825;
squeal_samples[39271]=6352;
squeal_samples[39272]=9165;
squeal_samples[39273]=11856;
squeal_samples[39274]=14430;
squeal_samples[39275]=16895;
squeal_samples[39276]=19242;
squeal_samples[39277]=21488;
squeal_samples[39278]=23637;
squeal_samples[39279]=25691;
squeal_samples[39280]=27647;
squeal_samples[39281]=29528;
squeal_samples[39282]=31310;
squeal_samples[39283]=33027;
squeal_samples[39284]=34659;
squeal_samples[39285]=36217;
squeal_samples[39286]=37708;
squeal_samples[39287]=39130;
squeal_samples[39288]=40487;
squeal_samples[39289]=41782;
squeal_samples[39290]=43027;
squeal_samples[39291]=44207;
squeal_samples[39292]=45338;
squeal_samples[39293]=46416;
squeal_samples[39294]=47449;
squeal_samples[39295]=48430;
squeal_samples[39296]=49370;
squeal_samples[39297]=50265;
squeal_samples[39298]=51125;
squeal_samples[39299]=51943;
squeal_samples[39300]=52731;
squeal_samples[39301]=53471;
squeal_samples[39302]=54189;
squeal_samples[39303]=54817;
squeal_samples[39304]=51294;
squeal_samples[39305]=45449;
squeal_samples[39306]=39983;
squeal_samples[39307]=34863;
squeal_samples[39308]=30072;
squeal_samples[39309]=25590;
squeal_samples[39310]=21388;
squeal_samples[39311]=17469;
squeal_samples[39312]=13790;
squeal_samples[39313]=10356;
squeal_samples[39314]=7129;
squeal_samples[39315]=4172;
squeal_samples[39316]=4890;
squeal_samples[39317]=7775;
squeal_samples[39318]=10515;
squeal_samples[39319]=13158;
squeal_samples[39320]=15666;
squeal_samples[39321]=18072;
squeal_samples[39322]=20368;
squeal_samples[39323]=22573;
squeal_samples[39324]=24660;
squeal_samples[39325]=26676;
squeal_samples[39326]=28587;
squeal_samples[39327]=30422;
squeal_samples[39328]=32170;
squeal_samples[39329]=33841;
squeal_samples[39330]=35435;
squeal_samples[39331]=36962;
squeal_samples[39332]=38413;
squeal_samples[39333]=39810;
squeal_samples[39334]=41131;
squeal_samples[39335]=42404;
squeal_samples[39336]=43611;
squeal_samples[39337]=44769;
squeal_samples[39338]=45874;
squeal_samples[39339]=46928;
squeal_samples[39340]=47937;
squeal_samples[39341]=48898;
squeal_samples[39342]=49816;
squeal_samples[39343]=50689;
squeal_samples[39344]=51530;
squeal_samples[39345]=52327;
squeal_samples[39346]=53098;
squeal_samples[39347]=53819;
squeal_samples[39348]=54530;
squeal_samples[39349]=53858;
squeal_samples[39350]=48314;
squeal_samples[39351]=42661;
squeal_samples[39352]=37367;
squeal_samples[39353]=32419;
squeal_samples[39354]=27783;
squeal_samples[39355]=23448;
squeal_samples[39356]=19386;
squeal_samples[39357]=15587;
squeal_samples[39358]=12037;
squeal_samples[39359]=8703;
squeal_samples[39360]=5599;
squeal_samples[39361]=3808;
squeal_samples[39362]=6338;
squeal_samples[39363]=9150;
squeal_samples[39364]=11840;
squeal_samples[39365]=14417;
squeal_samples[39366]=16872;
squeal_samples[39367]=19224;
squeal_samples[39368]=21465;
squeal_samples[39369]=23620;
squeal_samples[39370]=25667;
squeal_samples[39371]=27636;
squeal_samples[39372]=29503;
squeal_samples[39373]=31300;
squeal_samples[39374]=33003;
squeal_samples[39375]=34641;
squeal_samples[39376]=36194;
squeal_samples[39377]=37690;
squeal_samples[39378]=39108;
squeal_samples[39379]=40469;
squeal_samples[39380]=41764;
squeal_samples[39381]=43009;
squeal_samples[39382]=44184;
squeal_samples[39383]=45320;
squeal_samples[39384]=46395;
squeal_samples[39385]=47428;
squeal_samples[39386]=48410;
squeal_samples[39387]=49349;
squeal_samples[39388]=50252;
squeal_samples[39389]=51103;
squeal_samples[39390]=51925;
squeal_samples[39391]=52707;
squeal_samples[39392]=53453;
squeal_samples[39393]=54169;
squeal_samples[39394]=54802;
squeal_samples[39395]=51272;
squeal_samples[39396]=45431;
squeal_samples[39397]=39960;
squeal_samples[39398]=34845;
squeal_samples[39399]=30056;
squeal_samples[39400]=25569;
squeal_samples[39401]=21375;
squeal_samples[39402]=17446;
squeal_samples[39403]=13772;
squeal_samples[39404]=10334;
squeal_samples[39405]=7110;
squeal_samples[39406]=4150;
squeal_samples[39407]=4872;
squeal_samples[39408]=7751;
squeal_samples[39409]=10499;
squeal_samples[39410]=13135;
squeal_samples[39411]=15646;
squeal_samples[39412]=18052;
squeal_samples[39413]=20346;
squeal_samples[39414]=22554;
squeal_samples[39415]=24646;
squeal_samples[39416]=26654;
squeal_samples[39417]=28566;
squeal_samples[39418]=30403;
squeal_samples[39419]=32149;
squeal_samples[39420]=33821;
squeal_samples[39421]=35415;
squeal_samples[39422]=36939;
squeal_samples[39423]=38395;
squeal_samples[39424]=39789;
squeal_samples[39425]=41112;
squeal_samples[39426]=42382;
squeal_samples[39427]=43592;
squeal_samples[39428]=44745;
squeal_samples[39429]=45859;
squeal_samples[39430]=46903;
squeal_samples[39431]=47921;
squeal_samples[39432]=48874;
squeal_samples[39433]=49798;
squeal_samples[39434]=50668;
squeal_samples[39435]=51513;
squeal_samples[39436]=52311;
squeal_samples[39437]=53073;
squeal_samples[39438]=53803;
squeal_samples[39439]=54507;
squeal_samples[39440]=53838;
squeal_samples[39441]=48294;
squeal_samples[39442]=42640;
squeal_samples[39443]=37348;
squeal_samples[39444]=32398;
squeal_samples[39445]=27762;
squeal_samples[39446]=23430;
squeal_samples[39447]=19361;
squeal_samples[39448]=15572;
squeal_samples[39449]=12011;
squeal_samples[39450]=8689;
squeal_samples[39451]=5573;
squeal_samples[39452]=3793;
squeal_samples[39453]=6312;
squeal_samples[39454]=9134;
squeal_samples[39455]=11817;
squeal_samples[39456]=14398;
squeal_samples[39457]=16852;
squeal_samples[39458]=19203;
squeal_samples[39459]=21446;
squeal_samples[39460]=23597;
squeal_samples[39461]=25650;
squeal_samples[39462]=27612;
squeal_samples[39463]=29487;
squeal_samples[39464]=31275;
squeal_samples[39465]=32986;
squeal_samples[39466]=34619;
squeal_samples[39467]=36175;
squeal_samples[39468]=37670;
squeal_samples[39469]=39085;
squeal_samples[39470]=40450;
squeal_samples[39471]=41744;
squeal_samples[39472]=42988;
squeal_samples[39473]=44166;
squeal_samples[39474]=45296;
squeal_samples[39475]=46377;
squeal_samples[39476]=47407;
squeal_samples[39477]=48390;
squeal_samples[39478]=49329;
squeal_samples[39479]=50230;
squeal_samples[39480]=51085;
squeal_samples[39481]=51902;
squeal_samples[39482]=52689;
squeal_samples[39483]=53433;
squeal_samples[39484]=54146;
squeal_samples[39485]=54784;
squeal_samples[39486]=51252;
squeal_samples[39487]=45407;
squeal_samples[39488]=39946;
squeal_samples[39489]=34819;
squeal_samples[39490]=30038;
squeal_samples[39491]=25550;
squeal_samples[39492]=21351;
squeal_samples[39493]=17430;
squeal_samples[39494]=13748;
squeal_samples[39495]=10315;
squeal_samples[39496]=7091;
squeal_samples[39497]=4128;
squeal_samples[39498]=4853;
squeal_samples[39499]=7729;
squeal_samples[39500]=10479;
squeal_samples[39501]=13115;
squeal_samples[39502]=15628;
squeal_samples[39503]=18028;
squeal_samples[39504]=20330;
squeal_samples[39505]=22529;
squeal_samples[39506]=24628;
squeal_samples[39507]=26633;
squeal_samples[39508]=28548;
squeal_samples[39509]=30380;
squeal_samples[39510]=32131;
squeal_samples[39511]=33797;
squeal_samples[39512]=35398;
squeal_samples[39513]=36918;
squeal_samples[39514]=38374;
squeal_samples[39515]=39769;
squeal_samples[39516]=41090;
squeal_samples[39517]=42364;
squeal_samples[39518]=43570;
squeal_samples[39519]=44728;
squeal_samples[39520]=45834;
squeal_samples[39521]=46886;
squeal_samples[39522]=47897;
squeal_samples[39523]=48859;
squeal_samples[39524]=49772;
squeal_samples[39525]=50654;
squeal_samples[39526]=51486;
squeal_samples[39527]=52297;
squeal_samples[39528]=53047;
squeal_samples[39529]=53787;
squeal_samples[39530]=54484;
squeal_samples[39531]=53819;
squeal_samples[39532]=48274;
squeal_samples[39533]=42619;
squeal_samples[39534]=37328;
squeal_samples[39535]=32377;
squeal_samples[39536]=27743;
squeal_samples[39537]=23407;
squeal_samples[39538]=19345;
squeal_samples[39539]=15547;
squeal_samples[39540]=11995;
squeal_samples[39541]=8664;
squeal_samples[39542]=5557;
squeal_samples[39543]=3768;
squeal_samples[39544]=6297;
squeal_samples[39545]=9108;
squeal_samples[39546]=11803;
squeal_samples[39547]=14371;
squeal_samples[39548]=16838;
squeal_samples[39549]=19176;
squeal_samples[39550]=21431;
squeal_samples[39551]=23574;
squeal_samples[39552]=25631;
squeal_samples[39553]=27591;
squeal_samples[39554]=29466;
squeal_samples[39555]=31255;
squeal_samples[39556]=32966;
squeal_samples[39557]=34599;
squeal_samples[39558]=36154;
squeal_samples[39559]=37648;
squeal_samples[39560]=39069;
squeal_samples[39561]=40425;
squeal_samples[39562]=41728;
squeal_samples[39563]=42964;
squeal_samples[39564]=44147;
squeal_samples[39565]=45276;
squeal_samples[39566]=46356;
squeal_samples[39567]=47387;
squeal_samples[39568]=48369;
squeal_samples[39569]=49309;
squeal_samples[39570]=50209;
squeal_samples[39571]=51064;
squeal_samples[39572]=51882;
squeal_samples[39573]=52668;
squeal_samples[39574]=53411;
squeal_samples[39575]=54127;
squeal_samples[39576]=54810;
squeal_samples[39577]=52069;
squeal_samples[39578]=46170;
squeal_samples[39579]=40655;
squeal_samples[39580]=35486;
squeal_samples[39581]=30658;
squeal_samples[39582]=26125;
squeal_samples[39583]=21893;
squeal_samples[39584]=17931;
squeal_samples[39585]=14227;
squeal_samples[39586]=10753;
squeal_samples[39587]=7506;
squeal_samples[39588]=4462;
squeal_samples[39589]=4498;
squeal_samples[39590]=7391;
squeal_samples[39591]=10152;
squeal_samples[39592]=12802;
squeal_samples[39593]=15329;
squeal_samples[39594]=17749;
squeal_samples[39595]=20053;
squeal_samples[39596]=22266;
squeal_samples[39597]=24373;
squeal_samples[39598]=26390;
squeal_samples[39599]=28316;
squeal_samples[39600]=30159;
squeal_samples[39601]=31920;
squeal_samples[39602]=33594;
squeal_samples[39603]=35202;
squeal_samples[39604]=36730;
squeal_samples[39605]=38197;
squeal_samples[39606]=39590;
squeal_samples[39607]=40925;
squeal_samples[39608]=42200;
squeal_samples[39609]=43421;
squeal_samples[39610]=44581;
squeal_samples[39611]=45690;
squeal_samples[39612]=46752;
squeal_samples[39613]=47762;
squeal_samples[39614]=48728;
squeal_samples[39615]=49652;
squeal_samples[39616]=50530;
squeal_samples[39617]=51375;
squeal_samples[39618]=52176;
squeal_samples[39619]=52951;
squeal_samples[39620]=53685;
squeal_samples[39621]=54384;
squeal_samples[39622]=54574;
squeal_samples[39623]=49807;
squeal_samples[39624]=44061;
squeal_samples[39625]=38674;
squeal_samples[39626]=33640;
squeal_samples[39627]=28916;
squeal_samples[39628]=24506;
squeal_samples[39629]=20371;
squeal_samples[39630]=16507;
squeal_samples[39631]=12888;
squeal_samples[39632]=9501;
squeal_samples[39633]=6332;
squeal_samples[39634]=3777;
squeal_samples[39635]=5589;
squeal_samples[39636]=8433;
squeal_samples[39637]=11154;
squeal_samples[39638]=13758;
squeal_samples[39639]=16242;
squeal_samples[39640]=18618;
squeal_samples[39641]=20885;
squeal_samples[39642]=23058;
squeal_samples[39643]=25136;
squeal_samples[39644]=27115;
squeal_samples[39645]=29013;
squeal_samples[39646]=30816;
squeal_samples[39647]=32550;
squeal_samples[39648]=34197;
squeal_samples[39649]=35778;
squeal_samples[39650]=37278;
squeal_samples[39651]=38721;
squeal_samples[39652]=40086;
squeal_samples[39653]=41406;
squeal_samples[39654]=42655;
squeal_samples[39655]=43851;
squeal_samples[39656]=44995;
squeal_samples[39657]=46086;
squeal_samples[39658]=47127;
squeal_samples[39659]=48121;
squeal_samples[39660]=49072;
squeal_samples[39661]=49976;
squeal_samples[39662]=50850;
squeal_samples[39663]=51670;
squeal_samples[39664]=52463;
squeal_samples[39665]=53216;
squeal_samples[39666]=53944;
squeal_samples[39667]=54630;
squeal_samples[39668]=53374;
squeal_samples[39669]=47597;
squeal_samples[39670]=41985;
squeal_samples[39671]=36733;
squeal_samples[39672]=31819;
squeal_samples[39673]=27220;
squeal_samples[39674]=22913;
squeal_samples[39675]=18880;
squeal_samples[39676]=15111;
squeal_samples[39677]=11581;
squeal_samples[39678]=8280;
squeal_samples[39679]=5190;
squeal_samples[39680]=3925;
squeal_samples[39681]=6661;
squeal_samples[39682]=9461;
squeal_samples[39683]=12132;
squeal_samples[39684]=14694;
squeal_samples[39685]=17132;
squeal_samples[39686]=19472;
squeal_samples[39687]=21700;
squeal_samples[39688]=23839;
squeal_samples[39689]=25881;
squeal_samples[39690]=27827;
squeal_samples[39691]=29691;
squeal_samples[39692]=31463;
squeal_samples[39693]=33164;
squeal_samples[39694]=34788;
squeal_samples[39695]=36339;
squeal_samples[39696]=37815;
squeal_samples[39697]=39230;
squeal_samples[39698]=40578;
squeal_samples[39699]=41872;
squeal_samples[39700]=43100;
squeal_samples[39701]=44276;
squeal_samples[39702]=45396;
squeal_samples[39703]=46472;
squeal_samples[39704]=47492;
squeal_samples[39705]=48475;
squeal_samples[39706]=49408;
squeal_samples[39707]=50299;
squeal_samples[39708]=51152;
squeal_samples[39709]=51961;
squeal_samples[39710]=52741;
squeal_samples[39711]=53483;
squeal_samples[39712]=54197;
squeal_samples[39713]=54816;
squeal_samples[39714]=51289;
squeal_samples[39715]=45441;
squeal_samples[39716]=39963;
squeal_samples[39717]=34847;
squeal_samples[39718]=30047;
squeal_samples[39719]=25561;
squeal_samples[39720]=21354;
squeal_samples[39721]=17433;
squeal_samples[39722]=13746;
squeal_samples[39723]=10313;
squeal_samples[39724]=7083;
squeal_samples[39725]=4116;
squeal_samples[39726]=4839;
squeal_samples[39727]=7718;
squeal_samples[39728]=10464;
squeal_samples[39729]=13098;
squeal_samples[39730]=15608;
squeal_samples[39731]=18010;
squeal_samples[39732]=20308;
squeal_samples[39733]=22503;
squeal_samples[39734]=24607;
squeal_samples[39735]=26608;
squeal_samples[39736]=28522;
squeal_samples[39737]=30355;
squeal_samples[39738]=32103;
squeal_samples[39739]=33772;
squeal_samples[39740]=35366;
squeal_samples[39741]=36890;
squeal_samples[39742]=38346;
squeal_samples[39743]=39732;
squeal_samples[39744]=41064;
squeal_samples[39745]=42325;
squeal_samples[39746]=43539;
squeal_samples[39747]=44691;
squeal_samples[39748]=45796;
squeal_samples[39749]=46850;
squeal_samples[39750]=47859;
squeal_samples[39751]=48815;
squeal_samples[39752]=49737;
squeal_samples[39753]=50607;
squeal_samples[39754]=51454;
squeal_samples[39755]=52248;
squeal_samples[39756]=53015;
squeal_samples[39757]=53741;
squeal_samples[39758]=54440;
squeal_samples[39759]=54257;
squeal_samples[39760]=49037;
squeal_samples[39761]=43334;
squeal_samples[39762]=37996;
squeal_samples[39763]=32997;
squeal_samples[39764]=28318;
squeal_samples[39765]=23943;
squeal_samples[39766]=19840;
squeal_samples[39767]=16016;
squeal_samples[39768]=12423;
squeal_samples[39769]=9062;
squeal_samples[39770]=5923;
squeal_samples[39771]=3708;
squeal_samples[39772]=5923;
squeal_samples[39773]=8749;
squeal_samples[39774]=11456;
squeal_samples[39775]=14041;
squeal_samples[39776]=16518;
squeal_samples[39777]=18874;
squeal_samples[39778]=21131;
squeal_samples[39779]=23295;
squeal_samples[39780]=25352;
squeal_samples[39781]=27329;
squeal_samples[39782]=29204;
squeal_samples[39783]=31013;
squeal_samples[39784]=32729;
squeal_samples[39785]=34368;
squeal_samples[39786]=35937;
squeal_samples[39787]=37434;
squeal_samples[39788]=38860;
squeal_samples[39789]=40229;
squeal_samples[39790]=41530;
squeal_samples[39791]=42777;
squeal_samples[39792]=43968;
squeal_samples[39793]=45099;
squeal_samples[39794]=46186;
squeal_samples[39795]=47222;
squeal_samples[39796]=48211;
squeal_samples[39797]=49153;
squeal_samples[39798]=50058;
squeal_samples[39799]=50918;
squeal_samples[39800]=51747;
squeal_samples[39801]=52528;
squeal_samples[39802]=53281;
squeal_samples[39803]=53998;
squeal_samples[39804]=54689;
squeal_samples[39805]=52734;
squeal_samples[39806]=46844;
squeal_samples[39807]=41282;
squeal_samples[39808]=36073;
squeal_samples[39809]=31196;
squeal_samples[39810]=26635;
squeal_samples[39811]=22362;
squeal_samples[39812]=18367;
squeal_samples[39813]=14629;
squeal_samples[39814]=11128;
squeal_samples[39815]=7851;
squeal_samples[39816]=4786;
squeal_samples[39817]=4128;
squeal_samples[39818]=6990;
squeal_samples[39819]=9768;
squeal_samples[39820]=12426;
squeal_samples[39821]=14974;
squeal_samples[39822]=17401;
squeal_samples[39823]=19723;
squeal_samples[39824]=21947;
squeal_samples[39825]=24068;
squeal_samples[39826]=26096;
squeal_samples[39827]=28030;
squeal_samples[39828]=29884;
squeal_samples[39829]=31648;
squeal_samples[39830]=33346;
squeal_samples[39831]=34953;
squeal_samples[39832]=36498;
squeal_samples[39833]=37966;
squeal_samples[39834]=39370;
squeal_samples[39835]=40720;
squeal_samples[39836]=41995;
squeal_samples[39837]=43220;
squeal_samples[39838]=44389;
squeal_samples[39839]=45503;
squeal_samples[39840]=46572;
squeal_samples[39841]=47587;
squeal_samples[39842]=48563;
squeal_samples[39843]=49492;
squeal_samples[39844]=50378;
squeal_samples[39845]=51224;
squeal_samples[39846]=52035;
squeal_samples[39847]=52807;
squeal_samples[39848]=53542;
squeal_samples[39849]=54250;
squeal_samples[39850]=54716;
squeal_samples[39851]=50497;
squeal_samples[39852]=44709;
squeal_samples[39853]=39273;
squeal_samples[39854]=34199;
squeal_samples[39855]=29441;
squeal_samples[39856]=24993;
squeal_samples[39857]=20819;
squeal_samples[39858]=16929;
squeal_samples[39859]=13278;
squeal_samples[39860]=9864;
squeal_samples[39861]=6666;
squeal_samples[39862]=3863;
squeal_samples[39863]=5173;
squeal_samples[39864]=8035;
squeal_samples[39865]=10773;
squeal_samples[39866]=13385;
squeal_samples[39867]=15889;
squeal_samples[39868]=18273;
squeal_samples[39869]=20558;
squeal_samples[39870]=22742;
squeal_samples[39871]=24828;
squeal_samples[39872]=26825;
squeal_samples[39873]=28723;
squeal_samples[39874]=30548;
squeal_samples[39875]=32285;
squeal_samples[39876]=33947;
squeal_samples[39877]=35531;
squeal_samples[39878]=37045;
squeal_samples[39879]=38493;
squeal_samples[39880]=39872;
squeal_samples[39881]=41190;
squeal_samples[39882]=42453;
squeal_samples[39883]=43654;
squeal_samples[39884]=44803;
squeal_samples[39885]=45900;
squeal_samples[39886]=46947;
squeal_samples[39887]=47950;
squeal_samples[39888]=48908;
squeal_samples[39889]=49816;
squeal_samples[39890]=50691;
squeal_samples[39891]=51516;
squeal_samples[39892]=52322;
squeal_samples[39893]=53070;
squeal_samples[39894]=53808;
squeal_samples[39895]=54496;
squeal_samples[39896]=53824;
squeal_samples[39897]=48275;
squeal_samples[39898]=42618;
squeal_samples[39899]=37324;
squeal_samples[39900]=32366;
squeal_samples[39901]=27727;
squeal_samples[39902]=23386;
squeal_samples[39903]=19316;
squeal_samples[39904]=15524;
squeal_samples[39905]=11959;
squeal_samples[39906]=8629;
squeal_samples[39907]=5518;
squeal_samples[39908]=3725;
squeal_samples[39909]=6253;
squeal_samples[39910]=9067;
squeal_samples[39911]=11757;
squeal_samples[39912]=14326;
squeal_samples[39913]=16785;
squeal_samples[39914]=19132;
squeal_samples[39915]=21379;
squeal_samples[39916]=23521;
squeal_samples[39917]=25578;
squeal_samples[39918]=27535;
squeal_samples[39919]=29415;
squeal_samples[39920]=31193;
squeal_samples[39921]=32909;
squeal_samples[39922]=34535;
squeal_samples[39923]=36100;
squeal_samples[39924]=37585;
squeal_samples[39925]=39012;
squeal_samples[39926]=40364;
squeal_samples[39927]=41664;
squeal_samples[39928]=42898;
squeal_samples[39929]=44084;
squeal_samples[39930]=45210;
squeal_samples[39931]=46291;
squeal_samples[39932]=47317;
squeal_samples[39933]=48304;
squeal_samples[39934]=49245;
squeal_samples[39935]=50138;
squeal_samples[39936]=50993;
squeal_samples[39937]=51813;
squeal_samples[39938]=52596;
squeal_samples[39939]=53342;
squeal_samples[39940]=54055;
squeal_samples[39941]=54740;
squeal_samples[39942]=52785;
squeal_samples[39943]=46891;
squeal_samples[39944]=41319;
squeal_samples[39945]=36110;
squeal_samples[39946]=31223;
squeal_samples[39947]=26663;
squeal_samples[39948]=22383;
squeal_samples[39949]=18387;
squeal_samples[39950]=14641;
squeal_samples[39951]=11141;
squeal_samples[39952]=7865;
squeal_samples[39953]=4793;
squeal_samples[39954]=4132;
squeal_samples[39955]=6990;
squeal_samples[39956]=9770;
squeal_samples[39957]=12431;
squeal_samples[39958]=14972;
squeal_samples[39959]=17402;
squeal_samples[39960]=19717;
squeal_samples[39961]=21938;
squeal_samples[39962]=24063;
squeal_samples[39963]=26088;
squeal_samples[39964]=28031;
squeal_samples[39965]=29877;
squeal_samples[39966]=31643;
squeal_samples[39967]=33328;
squeal_samples[39968]=34944;
squeal_samples[39969]=36479;
squeal_samples[39970]=37955;
squeal_samples[39971]=39355;
squeal_samples[39972]=40699;
squeal_samples[39973]=41983;
squeal_samples[39974]=43204;
squeal_samples[39975]=44371;
squeal_samples[39976]=45488;
squeal_samples[39977]=46552;
squeal_samples[39978]=47574;
squeal_samples[39979]=48541;
squeal_samples[39980]=49476;
squeal_samples[39981]=50354;
squeal_samples[39982]=51208;
squeal_samples[39983]=52009;
squeal_samples[39984]=52780;
squeal_samples[39985]=53524;
squeal_samples[39986]=54224;
squeal_samples[39987]=54851;
squeal_samples[39988]=51309;
squeal_samples[39989]=45460;
squeal_samples[39990]=39981;
squeal_samples[39991]=34854;
squeal_samples[39992]=30054;
squeal_samples[39993]=25558;
squeal_samples[39994]=21355;
squeal_samples[39995]=17424;
squeal_samples[39996]=13742;
squeal_samples[39997]=10295;
squeal_samples[39998]=7071;
squeal_samples[39999]=4098;
squeal_samples[40000]=4818;
squeal_samples[40001]=7693;
squeal_samples[40002]=10439;
squeal_samples[40003]=13066;
squeal_samples[40004]=15583;
squeal_samples[40005]=17981;
squeal_samples[40006]=20279;
squeal_samples[40007]=22471;
squeal_samples[40008]=24573;
squeal_samples[40009]=26572;
squeal_samples[40010]=28494;
squeal_samples[40011]=30315;
squeal_samples[40012]=32070;
squeal_samples[40013]=33729;
squeal_samples[40014]=35329;
squeal_samples[40015]=36850;
squeal_samples[40016]=38307;
squeal_samples[40017]=39689;
squeal_samples[40018]=41017;
squeal_samples[40019]=42285;
squeal_samples[40020]=43489;
squeal_samples[40021]=44652;
squeal_samples[40022]=45746;
squeal_samples[40023]=46805;
squeal_samples[40024]=47806;
squeal_samples[40025]=48766;
squeal_samples[40026]=49688;
squeal_samples[40027]=50561;
squeal_samples[40028]=51405;
squeal_samples[40029]=52198;
squeal_samples[40030]=52964;
squeal_samples[40031]=53690;
squeal_samples[40032]=54393;
squeal_samples[40033]=54572;
squeal_samples[40034]=49805;
squeal_samples[40035]=44044;
squeal_samples[40036]=38656;
squeal_samples[40037]=33612;
squeal_samples[40038]=28891;
squeal_samples[40039]=24474;
squeal_samples[40040]=20333;
squeal_samples[40041]=16473;
squeal_samples[40042]=12844;
squeal_samples[40043]=9459;
squeal_samples[40044]=6285;
squeal_samples[40045]=3728;
squeal_samples[40046]=5543;
squeal_samples[40047]=8379;
squeal_samples[40048]=11096;
squeal_samples[40049]=13698;
squeal_samples[40050]=16186;
squeal_samples[40051]=18553;
squeal_samples[40052]=20826;
squeal_samples[40053]=23000;
squeal_samples[40054]=25071;
squeal_samples[40055]=27054;
squeal_samples[40056]=28941;
squeal_samples[40057]=30753;
squeal_samples[40058]=32480;
squeal_samples[40059]=34129;
squeal_samples[40060]=35702;
squeal_samples[40061]=37211;
squeal_samples[40062]=38646;
squeal_samples[40063]=40025;
squeal_samples[40064]=41323;
squeal_samples[40065]=42588;
squeal_samples[40066]=43770;
squeal_samples[40067]=44924;
squeal_samples[40068]=46003;
squeal_samples[40069]=47049;
squeal_samples[40070]=48040;
squeal_samples[40071]=48991;
squeal_samples[40072]=49898;
squeal_samples[40073]=50766;
squeal_samples[40074]=51593;
squeal_samples[40075]=52381;
squeal_samples[40076]=53136;
squeal_samples[40077]=53862;
squeal_samples[40078]=54551;
squeal_samples[40079]=53873;
squeal_samples[40080]=48319;
squeal_samples[40081]=42651;
squeal_samples[40082]=37356;
squeal_samples[40083]=32393;
squeal_samples[40084]=27751;
squeal_samples[40085]=23400;
squeal_samples[40086]=19341;
squeal_samples[40087]=15527;
squeal_samples[40088]=11970;
squeal_samples[40089]=8634;
squeal_samples[40090]=5511;
squeal_samples[40091]=3733;
squeal_samples[40092]=6246;
squeal_samples[40093]=9062;
squeal_samples[40094]=11748;
squeal_samples[40095]=14320;
squeal_samples[40096]=16776;
squeal_samples[40097]=19124;
squeal_samples[40098]=21365;
squeal_samples[40099]=23516;
squeal_samples[40100]=25562;
squeal_samples[40101]=27519;
squeal_samples[40102]=29394;
squeal_samples[40103]=31182;
squeal_samples[40104]=32888;
squeal_samples[40105]=34520;
squeal_samples[40106]=36077;
squeal_samples[40107]=37565;
squeal_samples[40108]=38985;
squeal_samples[40109]=40341;
squeal_samples[40110]=41641;
squeal_samples[40111]=42872;
squeal_samples[40112]=44061;
squeal_samples[40113]=45186;
squeal_samples[40114]=46261;
squeal_samples[40115]=47294;
squeal_samples[40116]=48273;
squeal_samples[40117]=49216;
squeal_samples[40118]=50109;
squeal_samples[40119]=50963;
squeal_samples[40120]=51784;
squeal_samples[40121]=52566;
squeal_samples[40122]=53313;
squeal_samples[40123]=54026;
squeal_samples[40124]=54709;
squeal_samples[40125]=52752;
squeal_samples[40126]=46854;
squeal_samples[40127]=41287;
squeal_samples[40128]=36073;
squeal_samples[40129]=31195;
squeal_samples[40130]=26627;
squeal_samples[40131]=22349;
squeal_samples[40132]=18351;
squeal_samples[40133]=14608;
squeal_samples[40134]=11104;
squeal_samples[40135]=7827;
squeal_samples[40136]=4756;
squeal_samples[40137]=4098;
squeal_samples[40138]=6956;
squeal_samples[40139]=9734;
squeal_samples[40140]=12392;
squeal_samples[40141]=14931;
squeal_samples[40142]=17367;
squeal_samples[40143]=19682;
squeal_samples[40144]=21905;
squeal_samples[40145]=24026;
squeal_samples[40146]=26050;
squeal_samples[40147]=27989;
squeal_samples[40148]=29837;
squeal_samples[40149]=31607;
squeal_samples[40150]=33297;
squeal_samples[40151]=34904;
squeal_samples[40152]=36449;
squeal_samples[40153]=37916;
squeal_samples[40154]=39323;
squeal_samples[40155]=40662;
squeal_samples[40156]=41945;
squeal_samples[40157]=43162;
squeal_samples[40158]=44337;
squeal_samples[40159]=45447;
squeal_samples[40160]=46514;
squeal_samples[40161]=47529;
squeal_samples[40162]=48508;
squeal_samples[40163]=49428;
squeal_samples[40164]=50320;
squeal_samples[40165]=51164;
squeal_samples[40166]=51970;
squeal_samples[40167]=52741;
squeal_samples[40168]=53482;
squeal_samples[40169]=54191;
squeal_samples[40170]=54809;
squeal_samples[40171]=51276;
squeal_samples[40172]=45418;
squeal_samples[40173]=39944;
squeal_samples[40174]=34810;
squeal_samples[40175]=30016;
squeal_samples[40176]=25523;
squeal_samples[40177]=21313;
squeal_samples[40178]=17387;
squeal_samples[40179]=13699;
squeal_samples[40180]=10255;
squeal_samples[40181]=7032;
squeal_samples[40182]=4056;
squeal_samples[40183]=4780;
squeal_samples[40184]=7650;
squeal_samples[40185]=10401;
squeal_samples[40186]=13024;
squeal_samples[40187]=15544;
squeal_samples[40188]=17941;
squeal_samples[40189]=20237;
squeal_samples[40190]=22434;
squeal_samples[40191]=24528;
squeal_samples[40192]=26538;
squeal_samples[40193]=28447;
squeal_samples[40194]=30280;
squeal_samples[40195]=32027;
squeal_samples[40196]=33689;
squeal_samples[40197]=35291;
squeal_samples[40198]=36806;
squeal_samples[40199]=38271;
squeal_samples[40200]=39645;
squeal_samples[40201]=40981;
squeal_samples[40202]=42241;
squeal_samples[40203]=43452;
squeal_samples[40204]=44609;
squeal_samples[40205]=45709;
squeal_samples[40206]=46763;
squeal_samples[40207]=47766;
squeal_samples[40208]=48728;
squeal_samples[40209]=49643;
squeal_samples[40210]=50527;
squeal_samples[40211]=51359;
squeal_samples[40212]=52163;
squeal_samples[40213]=52920;
squeal_samples[40214]=53653;
squeal_samples[40215]=54349;
squeal_samples[40216]=54535;
squeal_samples[40217]=49764;
squeal_samples[40218]=44003;
squeal_samples[40219]=38618;
squeal_samples[40220]=33569;
squeal_samples[40221]=28854;
squeal_samples[40222]=24431;
squeal_samples[40223]=20296;
squeal_samples[40224]=16429;
squeal_samples[40225]=12807;
squeal_samples[40226]=9417;
squeal_samples[40227]=6246;
squeal_samples[40228]=3688;
squeal_samples[40229]=5502;
squeal_samples[40230]=8339;
squeal_samples[40231]=11055;
squeal_samples[40232]=13660;
squeal_samples[40233]=16144;
squeal_samples[40234]=18513;
squeal_samples[40235]=20787;
squeal_samples[40236]=22958;
squeal_samples[40237]=25033;
squeal_samples[40238]=27012;
squeal_samples[40239]=28901;
squeal_samples[40240]=30714;
squeal_samples[40241]=32439;
squeal_samples[40242]=34088;
squeal_samples[40243]=35664;
squeal_samples[40244]=37168;
squeal_samples[40245]=38609;
squeal_samples[40246]=39980;
squeal_samples[40247]=41290;
squeal_samples[40248]=42539;
squeal_samples[40249]=43739;
squeal_samples[40250]=44875;
squeal_samples[40251]=45970;
squeal_samples[40252]=47004;
squeal_samples[40253]=48003;
squeal_samples[40254]=48949;
squeal_samples[40255]=49858;
squeal_samples[40256]=50727;
squeal_samples[40257]=51550;
squeal_samples[40258]=52343;
squeal_samples[40259]=53094;
squeal_samples[40260]=53823;
squeal_samples[40261]=54508;
squeal_samples[40262]=54314;
squeal_samples[40263]=49082;
squeal_samples[40264]=43378;
squeal_samples[40265]=38021;
squeal_samples[40266]=33021;
squeal_samples[40267]=28330;
squeal_samples[40268]=23945;
squeal_samples[40269]=19840;
squeal_samples[40270]=16000;
squeal_samples[40271]=12407;
squeal_samples[40272]=9042;
squeal_samples[40273]=5893;
squeal_samples[40274]=3673;
squeal_samples[40275]=5888;
squeal_samples[40276]=8711;
squeal_samples[40277]=11408;
squeal_samples[40278]=13997;
squeal_samples[40279]=16465;
squeal_samples[40280]=18824;
squeal_samples[40281]=21081;
squeal_samples[40282]=23235;
squeal_samples[40283]=25300;
squeal_samples[40284]=27262;
squeal_samples[40285]=29147;
squeal_samples[40286]=30943;
squeal_samples[40287]=32655;
squeal_samples[40288]=34303;
squeal_samples[40289]=35862;
squeal_samples[40290]=37362;
squeal_samples[40291]=38788;
squeal_samples[40292]=40149;
squeal_samples[40293]=41453;
squeal_samples[40294]=42698;
squeal_samples[40295]=43889;
squeal_samples[40296]=45021;
squeal_samples[40297]=46103;
squeal_samples[40298]=47138;
squeal_samples[40299]=48125;
squeal_samples[40300]=49072;
squeal_samples[40301]=49972;
squeal_samples[40302]=50828;
squeal_samples[40303]=51655;
squeal_samples[40304]=52435;
squeal_samples[40305]=53193;
squeal_samples[40306]=53903;
squeal_samples[40307]=54590;
squeal_samples[40308]=53914;
squeal_samples[40309]=48345;
squeal_samples[40310]=42682;
squeal_samples[40311]=37377;
squeal_samples[40312]=32413;
squeal_samples[40313]=27760;
squeal_samples[40314]=23416;
squeal_samples[40315]=19338;
squeal_samples[40316]=15537;
squeal_samples[40317]=11964;
squeal_samples[40318]=8635;
squeal_samples[40319]=5505;
squeal_samples[40320]=3719;
squeal_samples[40321]=6235;
squeal_samples[40322]=9050;
squeal_samples[40323]=11734;
squeal_samples[40324]=14309;
squeal_samples[40325]=16758;
squeal_samples[40326]=19102;
squeal_samples[40327]=21347;
squeal_samples[40328]=23492;
squeal_samples[40329]=25538;
squeal_samples[40330]=27498;
squeal_samples[40331]=29369;
squeal_samples[40332]=31156;
squeal_samples[40333]=32856;
squeal_samples[40334]=34494;
squeal_samples[40335]=36047;
squeal_samples[40336]=37537;
squeal_samples[40337]=38951;
squeal_samples[40338]=40308;
squeal_samples[40339]=41605;
squeal_samples[40340]=42840;
squeal_samples[40341]=44026;
squeal_samples[40342]=45146;
squeal_samples[40343]=46229;
squeal_samples[40344]=47252;
squeal_samples[40345]=48236;
squeal_samples[40346]=49175;
squeal_samples[40347]=50070;
squeal_samples[40348]=50923;
squeal_samples[40349]=51746;
squeal_samples[40350]=52519;
squeal_samples[40351]=53275;
squeal_samples[40352]=53979;
squeal_samples[40353]=54665;
squeal_samples[40354]=53396;
squeal_samples[40355]=47609;
squeal_samples[40356]=41990;
squeal_samples[40357]=36730;
squeal_samples[40358]=31802;
squeal_samples[40359]=27193;
squeal_samples[40360]=22877;
squeal_samples[40361]=18837;
squeal_samples[40362]=15063;
squeal_samples[40363]=11528;
squeal_samples[40364]=8219;
squeal_samples[40365]=5121;
squeal_samples[40366]=3851;
squeal_samples[40367]=6584;
squeal_samples[40368]=9382;
squeal_samples[40369]=12051;
squeal_samples[40370]=14606;
squeal_samples[40371]=17049;
squeal_samples[40372]=19378;
squeal_samples[40373]=21609;
squeal_samples[40374]=23743;
squeal_samples[40375]=25777;
squeal_samples[40376]=27727;
squeal_samples[40377]=29587;
squeal_samples[40378]=31362;
squeal_samples[40379]=33060;
squeal_samples[40380]=34677;
squeal_samples[40381]=36229;
squeal_samples[40382]=37704;
squeal_samples[40383]=39116;
squeal_samples[40384]=40465;
squeal_samples[40385]=41753;
squeal_samples[40386]=42983;
squeal_samples[40387]=44155;
squeal_samples[40388]=45280;
squeal_samples[40389]=46346;
squeal_samples[40390]=47370;
squeal_samples[40391]=48343;
squeal_samples[40392]=49280;
squeal_samples[40393]=50169;
squeal_samples[40394]=51021;
squeal_samples[40395]=51835;
squeal_samples[40396]=52605;
squeal_samples[40397]=53353;
squeal_samples[40398]=54057;
squeal_samples[40399]=54741;
squeal_samples[40400]=52780;
squeal_samples[40401]=46873;
squeal_samples[40402]=41304;
squeal_samples[40403]=36082;
squeal_samples[40404]=31202;
squeal_samples[40405]=26630;
squeal_samples[40406]=22349;
squeal_samples[40407]=18347;
squeal_samples[40408]=14598;
squeal_samples[40409]=11098;
squeal_samples[40410]=7810;
squeal_samples[40411]=4744;
squeal_samples[40412]=4072;
squeal_samples[40413]=6936;
squeal_samples[40414]=9712;
squeal_samples[40415]=12368;
squeal_samples[40416]=14911;
squeal_samples[40417]=17337;
squeal_samples[40418]=19650;
squeal_samples[40419]=21873;
squeal_samples[40420]=23991;
squeal_samples[40421]=26019;
squeal_samples[40422]=27954;
squeal_samples[40423]=29800;
squeal_samples[40424]=31569;
squeal_samples[40425]=33257;
squeal_samples[40426]=34866;
squeal_samples[40427]=36406;
squeal_samples[40428]=37870;
squeal_samples[40429]=39282;
squeal_samples[40430]=40617;
squeal_samples[40431]=41899;
squeal_samples[40432]=43122;
squeal_samples[40433]=44283;
squeal_samples[40434]=45408;
squeal_samples[40435]=46465;
squeal_samples[40436]=47485;
squeal_samples[40437]=48453;
squeal_samples[40438]=49383;
squeal_samples[40439]=50269;
squeal_samples[40440]=51115;
squeal_samples[40441]=51919;
squeal_samples[40442]=52694;
squeal_samples[40443]=53428;
squeal_samples[40444]=54141;
squeal_samples[40445]=54810;
squeal_samples[40446]=52058;
squeal_samples[40447]=46148;
squeal_samples[40448]=40623;
squeal_samples[40449]=35451;
squeal_samples[40450]=30602;
squeal_samples[40451]=26068;
squeal_samples[40452]=21823;
squeal_samples[40453]=17853;
squeal_samples[40454]=14133;
squeal_samples[40455]=10663;
squeal_samples[40456]=7404;
squeal_samples[40457]=4364;
squeal_samples[40458]=4389;
squeal_samples[40459]=7279;
squeal_samples[40460]=10038;
squeal_samples[40461]=12679;
squeal_samples[40462]=15212;
squeal_samples[40463]=17618;
squeal_samples[40464]=19931;
squeal_samples[40465]=22131;
squeal_samples[40466]=24238;
squeal_samples[40467]=26258;
squeal_samples[40468]=28178;
squeal_samples[40469]=30018;
squeal_samples[40470]=31770;
squeal_samples[40471]=33454;
squeal_samples[40472]=35051;
squeal_samples[40473]=36585;
squeal_samples[40474]=38042;
squeal_samples[40475]=39437;
squeal_samples[40476]=40771;
squeal_samples[40477]=42047;
squeal_samples[40478]=43263;
squeal_samples[40479]=44421;
squeal_samples[40480]=45533;
squeal_samples[40481]=46585;
squeal_samples[40482]=47600;
squeal_samples[40483]=48563;
squeal_samples[40484]=49487;
squeal_samples[40485]=50366;
squeal_samples[40486]=51209;
squeal_samples[40487]=52014;
squeal_samples[40488]=52778;
squeal_samples[40489]=53512;
squeal_samples[40490]=54211;
squeal_samples[40491]=54832;
squeal_samples[40492]=51286;
squeal_samples[40493]=45426;
squeal_samples[40494]=39947;
squeal_samples[40495]=34814;
squeal_samples[40496]=30008;
squeal_samples[40497]=25514;
squeal_samples[40498]=21302;
squeal_samples[40499]=17372;
squeal_samples[40500]=13676;
squeal_samples[40501]=10236;
squeal_samples[40502]=7004;
squeal_samples[40503]=4031;
squeal_samples[40504]=4751;
squeal_samples[40505]=7621;
squeal_samples[40506]=10364;
squeal_samples[40507]=12998;
squeal_samples[40508]=15502;
squeal_samples[40509]=17905;
squeal_samples[40510]=20196;
squeal_samples[40511]=22391;
squeal_samples[40512]=24491;
squeal_samples[40513]=26490;
squeal_samples[40514]=28403;
squeal_samples[40515]=30229;
squeal_samples[40516]=31979;
squeal_samples[40517]=33642;
squeal_samples[40518]=35239;
squeal_samples[40519]=36758;
squeal_samples[40520]=38211;
squeal_samples[40521]=39602;
squeal_samples[40522]=40923;
squeal_samples[40523]=42190;
squeal_samples[40524]=43396;
squeal_samples[40525]=44557;
squeal_samples[40526]=45653;
squeal_samples[40527]=46712;
squeal_samples[40528]=47709;
squeal_samples[40529]=48676;
squeal_samples[40530]=49584;
squeal_samples[40531]=50465;
squeal_samples[40532]=51304;
squeal_samples[40533]=52098;
squeal_samples[40534]=52866;
squeal_samples[40535]=53588;
squeal_samples[40536]=54295;
squeal_samples[40537]=54736;
squeal_samples[40538]=50529;
squeal_samples[40539]=44713;
squeal_samples[40540]=39276;
squeal_samples[40541]=34184;
squeal_samples[40542]=29423;
squeal_samples[40543]=24959;
squeal_samples[40544]=20786;
squeal_samples[40545]=16884;
squeal_samples[40546]=13227;
squeal_samples[40547]=9803;
squeal_samples[40548]=6604;
squeal_samples[40549]=3794;
squeal_samples[40550]=5104;
squeal_samples[40551]=7959;
squeal_samples[40552]=10694;
squeal_samples[40553]=13304;
squeal_samples[40554]=15805;
squeal_samples[40555]=18181;
squeal_samples[40556]=20468;
squeal_samples[40557]=22650;
squeal_samples[40558]=24732;
squeal_samples[40559]=26729;
squeal_samples[40560]=28621;
squeal_samples[40561]=30447;
squeal_samples[40562]=32175;
squeal_samples[40563]=33843;
squeal_samples[40564]=35421;
squeal_samples[40565]=36935;
squeal_samples[40566]=38378;
squeal_samples[40567]=39760;
squeal_samples[40568]=41078;
squeal_samples[40569]=42334;
squeal_samples[40570]=43537;
squeal_samples[40571]=44683;
squeal_samples[40572]=45778;
squeal_samples[40573]=46822;
squeal_samples[40574]=47823;
squeal_samples[40575]=48777;
squeal_samples[40576]=49688;
squeal_samples[40577]=50562;
squeal_samples[40578]=51385;
squeal_samples[40579]=52188;
squeal_samples[40580]=52942;
squeal_samples[40581]=53670;
squeal_samples[40582]=54363;
squeal_samples[40583]=54546;
squeal_samples[40584]=49765;
squeal_samples[40585]=44006;
squeal_samples[40586]=38611;
squeal_samples[40587]=33562;
squeal_samples[40588]=28837;
squeal_samples[40589]=24414;
squeal_samples[40590]=20272;
squeal_samples[40591]=16406;
squeal_samples[40592]=12773;
squeal_samples[40593]=9389;
squeal_samples[40594]=6207;
squeal_samples[40595]=3647;
squeal_samples[40596]=5460;
squeal_samples[40597]=8296;
squeal_samples[40598]=11016;
squeal_samples[40599]=13608;
squeal_samples[40600]=16100;
squeal_samples[40601]=18463;
squeal_samples[40602]=20736;
squeal_samples[40603]=22905;
squeal_samples[40604]=24978;
squeal_samples[40605]=26956;
squeal_samples[40606]=28846;
squeal_samples[40607]=30658;
squeal_samples[40608]=32378;
squeal_samples[40609]=34034;
squeal_samples[40610]=35599;
squeal_samples[40611]=37112;
squeal_samples[40612]=38539;
squeal_samples[40613]=39921;
squeal_samples[40614]=41222;
squeal_samples[40615]=42479;
squeal_samples[40616]=43671;
squeal_samples[40617]=44811;
squeal_samples[40618]=45901;
squeal_samples[40619]=46944;
squeal_samples[40620]=47936;
squeal_samples[40621]=48887;
squeal_samples[40622]=49788;
squeal_samples[40623]=50656;
squeal_samples[40624]=51485;
squeal_samples[40625]=52268;
squeal_samples[40626]=53030;
squeal_samples[40627]=53744;
squeal_samples[40628]=54440;
squeal_samples[40629]=54613;
squeal_samples[40630]=49829;
squeal_samples[40631]=44068;
squeal_samples[40632]=38665;
squeal_samples[40633]=33619;
squeal_samples[40634]=28884;
squeal_samples[40635]=24458;
squeal_samples[40636]=20313;
squeal_samples[40637]=16442;
squeal_samples[40638]=12810;
squeal_samples[40639]=9413;
squeal_samples[40640]=6236;
squeal_samples[40641]=3676;
squeal_samples[40642]=5481;
squeal_samples[40643]=8320;
squeal_samples[40644]=11036;
squeal_samples[40645]=13633;
squeal_samples[40646]=16116;
squeal_samples[40647]=18481;
squeal_samples[40648]=20752;
squeal_samples[40649]=22917;
squeal_samples[40650]=24990;
squeal_samples[40651]=26973;
squeal_samples[40652]=28858;
squeal_samples[40653]=30669;
squeal_samples[40654]=32391;
squeal_samples[40655]=34037;
squeal_samples[40656]=35615;
squeal_samples[40657]=37119;
squeal_samples[40658]=38550;
squeal_samples[40659]=39924;
squeal_samples[40660]=41229;
squeal_samples[40661]=42485;
squeal_samples[40662]=43678;
squeal_samples[40663]=44816;
squeal_samples[40664]=45903;
squeal_samples[40665]=46944;
squeal_samples[40666]=47938;
squeal_samples[40667]=48886;
squeal_samples[40668]=49791;
squeal_samples[40669]=50655;
squeal_samples[40670]=51486;
squeal_samples[40671]=52271;
squeal_samples[40672]=53026;
squeal_samples[40673]=53750;
squeal_samples[40674]=54432;
squeal_samples[40675]=54616;
squeal_samples[40676]=49824;
squeal_samples[40677]=44062;
squeal_samples[40678]=38661;
squeal_samples[40679]=33615;
squeal_samples[40680]=28879;
squeal_samples[40681]=24455;
squeal_samples[40682]=20306;
squeal_samples[40683]=16440;
squeal_samples[40684]=12802;
squeal_samples[40685]=9412;
squeal_samples[40686]=6230;
squeal_samples[40687]=3671;
squeal_samples[40688]=5477;
squeal_samples[40689]=8315;
squeal_samples[40690]=11027;
squeal_samples[40691]=13623;
squeal_samples[40692]=16109;
squeal_samples[40693]=18480;
squeal_samples[40694]=20744;
squeal_samples[40695]=22916;
squeal_samples[40696]=24977;
squeal_samples[40697]=26964;
squeal_samples[40698]=28848;
squeal_samples[40699]=30660;
squeal_samples[40700]=32379;
squeal_samples[40701]=34035;
squeal_samples[40702]=35602;
squeal_samples[40703]=37111;
squeal_samples[40704]=38540;
squeal_samples[40705]=39912;
squeal_samples[40706]=41223;
squeal_samples[40707]=42470;
squeal_samples[40708]=43673;
squeal_samples[40709]=44802;
squeal_samples[40710]=45902;
squeal_samples[40711]=46931;
squeal_samples[40712]=47929;
squeal_samples[40713]=48878;
squeal_samples[40714]=49783;
squeal_samples[40715]=50649;
squeal_samples[40716]=51473;
squeal_samples[40717]=52261;
squeal_samples[40718]=53020;
squeal_samples[40719]=53734;
squeal_samples[40720]=54428;
squeal_samples[40721]=54601;
squeal_samples[40722]=49818;
squeal_samples[40723]=44049;
squeal_samples[40724]=38655;
squeal_samples[40725]=33599;
squeal_samples[40726]=28875;
squeal_samples[40727]=24441;
squeal_samples[40728]=20298;
squeal_samples[40729]=16430;
squeal_samples[40730]=12791;
squeal_samples[40731]=9402;
squeal_samples[40732]=6221;
squeal_samples[40733]=3660;
squeal_samples[40734]=5468;
squeal_samples[40735]=8304;
squeal_samples[40736]=11017;
squeal_samples[40737]=13613;
squeal_samples[40738]=16100;
squeal_samples[40739]=18469;
squeal_samples[40740]=20734;
squeal_samples[40741]=22907;
squeal_samples[40742]=24965;
squeal_samples[40743]=26957;
squeal_samples[40744]=28836;
squeal_samples[40745]=30648;
squeal_samples[40746]=32374;
squeal_samples[40747]=34020;
squeal_samples[40748]=35598;
squeal_samples[40749]=37095;
squeal_samples[40750]=38533;
squeal_samples[40751]=39901;
squeal_samples[40752]=41214;
squeal_samples[40753]=42461;
squeal_samples[40754]=43659;
squeal_samples[40755]=44797;
squeal_samples[40756]=45887;
squeal_samples[40757]=46926;
squeal_samples[40758]=47916;
squeal_samples[40759]=48867;
squeal_samples[40760]=49776;
squeal_samples[40761]=50635;
squeal_samples[40762]=51467;
squeal_samples[40763]=52249;
squeal_samples[40764]=53010;
squeal_samples[40765]=53725;
squeal_samples[40766]=54416;
squeal_samples[40767]=54592;
squeal_samples[40768]=49808;
squeal_samples[40769]=44040;
squeal_samples[40770]=38643;
squeal_samples[40771]=33591;
squeal_samples[40772]=28864;
squeal_samples[40773]=24430;
squeal_samples[40774]=20291;
squeal_samples[40775]=16415;
squeal_samples[40776]=12786;
squeal_samples[40777]=9390;
squeal_samples[40778]=6211;
squeal_samples[40779]=3650;
squeal_samples[40780]=5457;
squeal_samples[40781]=8297;
squeal_samples[40782]=11004;
squeal_samples[40783]=13605;
squeal_samples[40784]=16089;
squeal_samples[40785]=18458;
squeal_samples[40786]=20727;
squeal_samples[40787]=22893;
squeal_samples[40788]=24959;
squeal_samples[40789]=26944;
squeal_samples[40790]=28827;
squeal_samples[40791]=30640;
squeal_samples[40792]=32360;
squeal_samples[40793]=34014;
squeal_samples[40794]=35584;
squeal_samples[40795]=37089;
squeal_samples[40796]=38521;
squeal_samples[40797]=39891;
squeal_samples[40798]=41204;
squeal_samples[40799]=42451;
squeal_samples[40800]=43650;
squeal_samples[40801]=44786;
squeal_samples[40802]=45877;
squeal_samples[40803]=46916;
squeal_samples[40804]=47905;
squeal_samples[40805]=48860;
squeal_samples[40806]=49763;
squeal_samples[40807]=50627;
squeal_samples[40808]=51456;
squeal_samples[40809]=52239;
squeal_samples[40810]=53000;
squeal_samples[40811]=53716;
squeal_samples[40812]=54404;
squeal_samples[40813]=54585;
squeal_samples[40814]=49794;
squeal_samples[40815]=44034;
squeal_samples[40816]=38630;
squeal_samples[40817]=33583;
squeal_samples[40818]=28853;
squeal_samples[40819]=24420;
squeal_samples[40820]=20281;
squeal_samples[40821]=16406;
squeal_samples[40822]=12775;
squeal_samples[40823]=9380;
squeal_samples[40824]=6202;
squeal_samples[40825]=3639;
squeal_samples[40826]=5448;
squeal_samples[40827]=8285;
squeal_samples[40828]=10996;
squeal_samples[40829]=13594;
squeal_samples[40830]=16080;
squeal_samples[40831]=18447;
squeal_samples[40832]=20718;
squeal_samples[40833]=22881;
squeal_samples[40834]=24952;
squeal_samples[40835]=26931;
squeal_samples[40836]=28820;
squeal_samples[40837]=30628;
squeal_samples[40838]=32350;
squeal_samples[40839]=34005;
squeal_samples[40840]=35573;
squeal_samples[40841]=37079;
squeal_samples[40842]=38512;
squeal_samples[40843]=39880;
squeal_samples[40844]=41194;
squeal_samples[40845]=42442;
squeal_samples[40846]=43638;
squeal_samples[40847]=44778;
squeal_samples[40848]=45866;
squeal_samples[40849]=46906;
squeal_samples[40850]=47896;
squeal_samples[40851]=48849;
squeal_samples[40852]=49753;
squeal_samples[40853]=50618;
squeal_samples[40854]=51445;
squeal_samples[40855]=52230;
squeal_samples[40856]=52989;
squeal_samples[40857]=53706;
squeal_samples[40858]=54396;
squeal_samples[40859]=54572;
squeal_samples[40860]=49788;
squeal_samples[40861]=44019;
squeal_samples[40862]=38624;
squeal_samples[40863]=33572;
squeal_samples[40864]=28841;
squeal_samples[40865]=24413;
squeal_samples[40866]=20269;
squeal_samples[40867]=16397;
squeal_samples[40868]=12765;
squeal_samples[40869]=9369;
squeal_samples[40870]=6192;
squeal_samples[40871]=3630;
squeal_samples[40872]=5437;
squeal_samples[40873]=8277;
squeal_samples[40874]=10983;
squeal_samples[40875]=13587;
squeal_samples[40876]=16066;
squeal_samples[40877]=18441;
squeal_samples[40878]=20705;
squeal_samples[40879]=22874;
squeal_samples[40880]=24939;
squeal_samples[40881]=26922;
squeal_samples[40882]=28811;
squeal_samples[40883]=30615;
squeal_samples[40884]=32345;
squeal_samples[40885]=33989;
squeal_samples[40886]=35567;
squeal_samples[40887]=37068;
squeal_samples[40888]=38501;
squeal_samples[40889]=39873;
squeal_samples[40890]=41180;
squeal_samples[40891]=42434;
squeal_samples[40892]=43628;
squeal_samples[40893]=44768;
squeal_samples[40894]=45856;
squeal_samples[40895]=46897;
squeal_samples[40896]=47883;
squeal_samples[40897]=48843;
squeal_samples[40898]=49740;
squeal_samples[40899]=50610;
squeal_samples[40900]=51433;
squeal_samples[40901]=52222;
squeal_samples[40902]=52977;
squeal_samples[40903]=53700;
squeal_samples[40904]=54380;
squeal_samples[40905]=54568;
squeal_samples[40906]=49772;
squeal_samples[40907]=44014;
squeal_samples[40908]=38611;
squeal_samples[40909]=33563;
squeal_samples[40910]=28832;
squeal_samples[40911]=24402;
squeal_samples[40912]=20258;
squeal_samples[40913]=16388;
squeal_samples[40914]=12754;
squeal_samples[40915]=9362;
squeal_samples[40916]=6179;
squeal_samples[40917]=3623;
squeal_samples[40918]=5423;
squeal_samples[40919]=8270;
squeal_samples[40920]=10972;
squeal_samples[40921]=13577;
squeal_samples[40922]=16057;
squeal_samples[40923]=18429;
squeal_samples[40924]=20697;
squeal_samples[40925]=22862;
squeal_samples[40926]=24930;
squeal_samples[40927]=26913;
squeal_samples[40928]=28798;
squeal_samples[40929]=30609;
squeal_samples[40930]=32331;
squeal_samples[40931]=33982;
squeal_samples[40932]=35555;
squeal_samples[40933]=37060;
squeal_samples[40934]=38488;
squeal_samples[40935]=39866;
squeal_samples[40936]=41168;
squeal_samples[40937]=42425;
squeal_samples[40938]=43617;
squeal_samples[40939]=44758;
squeal_samples[40940]=45847;
squeal_samples[40941]=46884;
squeal_samples[40942]=47877;
squeal_samples[40943]=48828;
squeal_samples[40944]=49733;
squeal_samples[40945]=50599;
squeal_samples[40946]=51422;
squeal_samples[40947]=52211;
squeal_samples[40948]=52970;
squeal_samples[40949]=53683;
squeal_samples[40950]=54377;
squeal_samples[40951]=54817;
squeal_samples[40952]=50593;
squeal_samples[40953]=44772;
squeal_samples[40954]=39324;
squeal_samples[40955]=34226;
squeal_samples[40956]=29451;
squeal_samples[40957]=24985;
squeal_samples[40958]=20801;
squeal_samples[40959]=16895;
squeal_samples[40960]=13230;
squeal_samples[40961]=9809;
squeal_samples[40962]=6592;
squeal_samples[40963]=3782;
squeal_samples[40964]=5083;
squeal_samples[40965]=7941;
squeal_samples[40966]=10666;
squeal_samples[40967]=13276;
squeal_samples[40968]=15772;
squeal_samples[40969]=18154;
squeal_samples[40970]=20428;
squeal_samples[40971]=22617;
squeal_samples[40972]=24690;
squeal_samples[40973]=26686;
squeal_samples[40974]=28583;
squeal_samples[40975]=30395;
squeal_samples[40976]=32135;
squeal_samples[40977]=33784;
squeal_samples[40978]=35375;
squeal_samples[40979]=36877;
squeal_samples[40980]=38325;
squeal_samples[40981]=39700;
squeal_samples[40982]=41021;
squeal_samples[40983]=42271;
squeal_samples[40984]=43479;
squeal_samples[40985]=44620;
squeal_samples[40986]=45715;
squeal_samples[40987]=46758;
squeal_samples[40988]=47761;
squeal_samples[40989]=48706;
squeal_samples[40990]=49623;
squeal_samples[40991]=50489;
squeal_samples[40992]=51319;
squeal_samples[40993]=52118;
squeal_samples[40994]=52866;
squeal_samples[40995]=53599;
squeal_samples[40996]=54284;
squeal_samples[40997]=54902;
squeal_samples[40998]=51342;
squeal_samples[40999]=45475;
squeal_samples[41000]=39982;
squeal_samples[41001]=34840;
squeal_samples[41002]=30028;
squeal_samples[41003]=25522;
squeal_samples[41004]=21303;
squeal_samples[41005]=17361;
squeal_samples[41006]=13668;
squeal_samples[41007]=10214;
squeal_samples[41008]=6983;
squeal_samples[41009]=3995;
squeal_samples[41010]=4718;
squeal_samples[41011]=7580;
squeal_samples[41012]=10327;
squeal_samples[41013]=12950;
squeal_samples[41014]=15458;
squeal_samples[41015]=17854;
squeal_samples[41016]=20145;
squeal_samples[41017]=22337;
squeal_samples[41018]=24434;
squeal_samples[41019]=26428;
squeal_samples[41020]=28342;
squeal_samples[41021]=30168;
squeal_samples[41022]=31911;
squeal_samples[41023]=33577;
squeal_samples[41024]=35165;
squeal_samples[41025]=36687;
squeal_samples[41026]=38138;
squeal_samples[41027]=39523;
squeal_samples[41028]=40848;
squeal_samples[41029]=42109;
squeal_samples[41030]=43322;
squeal_samples[41031]=44471;
squeal_samples[41032]=45571;
squeal_samples[41033]=46628;
squeal_samples[41034]=47625;
squeal_samples[41035]=48590;
squeal_samples[41036]=49497;
squeal_samples[41037]=50381;
squeal_samples[41038]=51209;
squeal_samples[41039]=52010;
squeal_samples[41040]=52764;
squeal_samples[41041]=53502;
squeal_samples[41042]=54190;
squeal_samples[41043]=54868;
squeal_samples[41044]=52089;
squeal_samples[41045]=46185;
squeal_samples[41046]=40637;
squeal_samples[41047]=35457;
squeal_samples[41048]=30603;
squeal_samples[41049]=26061;
squeal_samples[41050]=21809;
squeal_samples[41051]=17827;
squeal_samples[41052]=14111;
squeal_samples[41053]=10621;
squeal_samples[41054]=7364;
squeal_samples[41055]=4312;
squeal_samples[41056]=4337;
squeal_samples[41057]=7223;
squeal_samples[41058]=9980;
squeal_samples[41059]=12619;
squeal_samples[41060]=15144;
squeal_samples[41061]=17557;
squeal_samples[41062]=19857;
squeal_samples[41063]=22057;
squeal_samples[41064]=24161;
squeal_samples[41065]=26177;
squeal_samples[41066]=28095;
squeal_samples[41067]=29938;
squeal_samples[41068]=31689;
squeal_samples[41069]=33365;
squeal_samples[41070]=34962;
squeal_samples[41071]=36490;
squeal_samples[41072]=37950;
squeal_samples[41073]=39345;
squeal_samples[41074]=40674;
squeal_samples[41075]=41948;
squeal_samples[41076]=43160;
squeal_samples[41077]=44319;
squeal_samples[41078]=45427;
squeal_samples[41079]=46485;
squeal_samples[41080]=47493;
squeal_samples[41081]=48461;
squeal_samples[41082]=49379;
squeal_samples[41083]=50256;
squeal_samples[41084]=51102;
squeal_samples[41085]=51896;
squeal_samples[41086]=52667;
squeal_samples[41087]=53399;
squeal_samples[41088]=54099;
squeal_samples[41089]=54770;
squeal_samples[41090]=52800;
squeal_samples[41091]=46890;
squeal_samples[41092]=41302;
squeal_samples[41093]=36076;
squeal_samples[41094]=31180;
squeal_samples[41095]=26604;
squeal_samples[41096]=22315;
squeal_samples[41097]=18300;
squeal_samples[41098]=14552;
squeal_samples[41099]=11034;
squeal_samples[41100]=7751;
squeal_samples[41101]=4672;
squeal_samples[41102]=4005;
squeal_samples[41103]=6854;
squeal_samples[41104]=9634;
squeal_samples[41105]=12282;
squeal_samples[41106]=14826;
squeal_samples[41107]=17246;
squeal_samples[41108]=19562;
squeal_samples[41109]=21777;
squeal_samples[41110]=23901;
squeal_samples[41111]=25918;
squeal_samples[41112]=27855;
squeal_samples[41113]=29699;
squeal_samples[41114]=31460;
squeal_samples[41115]=33152;
squeal_samples[41116]=34753;
squeal_samples[41117]=36298;
squeal_samples[41118]=37760;
squeal_samples[41119]=39167;
squeal_samples[41120]=40501;
squeal_samples[41121]=41780;
squeal_samples[41122]=43004;
squeal_samples[41123]=44167;
squeal_samples[41124]=45282;
squeal_samples[41125]=46345;
squeal_samples[41126]=47359;
squeal_samples[41127]=48330;
squeal_samples[41128]=49255;
squeal_samples[41129]=50139;
squeal_samples[41130]=50986;
squeal_samples[41131]=51792;
squeal_samples[41132]=52561;
squeal_samples[41133]=53299;
squeal_samples[41134]=54005;
squeal_samples[41135]=54679;
squeal_samples[41136]=53398;
squeal_samples[41137]=47603;
squeal_samples[41138]=41971;
squeal_samples[41139]=36700;
squeal_samples[41140]=31768;
squeal_samples[41141]=27148;
squeal_samples[41142]=22825;
squeal_samples[41143]=18782;
squeal_samples[41144]=14993;
squeal_samples[41145]=11457;
squeal_samples[41146]=8136;
squeal_samples[41147]=5038;
squeal_samples[41148]=3761;
squeal_samples[41149]=6490;
squeal_samples[41150]=9282;
squeal_samples[41151]=11951;
squeal_samples[41152]=14502;
squeal_samples[41153]=16943;
squeal_samples[41154]=19267;
squeal_samples[41155]=21501;
squeal_samples[41156]=23623;
squeal_samples[41157]=25665;
squeal_samples[41158]=27601;
squeal_samples[41159]=29464;
squeal_samples[41160]=31233;
squeal_samples[41161]=32934;
squeal_samples[41162]=34550;
squeal_samples[41163]=36095;
squeal_samples[41164]=37574;
squeal_samples[41165]=38981;
squeal_samples[41166]=40330;
squeal_samples[41167]=41612;
squeal_samples[41168]=42842;
squeal_samples[41169]=44016;
squeal_samples[41170]=45137;
squeal_samples[41171]=46202;
squeal_samples[41172]=47226;
squeal_samples[41173]=48202;
squeal_samples[41174]=49134;
squeal_samples[41175]=50022;
squeal_samples[41176]=50871;
squeal_samples[41177]=51684;
squeal_samples[41178]=52460;
squeal_samples[41179]=53201;
squeal_samples[41180]=53908;
squeal_samples[41181]=54586;
squeal_samples[41182]=53895;
squeal_samples[41183]=48324;
squeal_samples[41184]=42648;
squeal_samples[41185]=37329;
squeal_samples[41186]=32357;
squeal_samples[41187]=27696;
squeal_samples[41188]=23337;
squeal_samples[41189]=19259;
squeal_samples[41190]=15448;
squeal_samples[41191]=11874;
squeal_samples[41192]=8527;
squeal_samples[41193]=5404;
squeal_samples[41194]=3609;
squeal_samples[41195]=6122;
squeal_samples[41196]=8929;
squeal_samples[41197]=11609;
squeal_samples[41198]=14183;
squeal_samples[41199]=16633;
squeal_samples[41200]=18978;
squeal_samples[41201]=21209;
squeal_samples[41202]=23358;
squeal_samples[41203]=25400;
squeal_samples[41204]=27358;
squeal_samples[41205]=29226;
squeal_samples[41206]=31010;
squeal_samples[41207]=32709;
squeal_samples[41208]=34342;
squeal_samples[41209]=35894;
squeal_samples[41210]=37385;
squeal_samples[41211]=38797;
squeal_samples[41212]=40158;
squeal_samples[41213]=41444;
squeal_samples[41214]=42686;
squeal_samples[41215]=43859;
squeal_samples[41216]=44991;
squeal_samples[41217]=46063;
squeal_samples[41218]=47091;
squeal_samples[41219]=48070;
squeal_samples[41220]=49007;
squeal_samples[41221]=49902;
squeal_samples[41222]=50758;
squeal_samples[41223]=51577;
squeal_samples[41224]=52350;
squeal_samples[41225]=53099;
squeal_samples[41226]=53811;
squeal_samples[41227]=54493;
squeal_samples[41228]=54287;
squeal_samples[41229]=49049;
squeal_samples[41230]=43319;
squeal_samples[41231]=37969;
squeal_samples[41232]=32946;
squeal_samples[41233]=28252;
squeal_samples[41234]=23861;
squeal_samples[41235]=19739;
squeal_samples[41236]=15903;
squeal_samples[41237]=12296;
squeal_samples[41238]=8927;
squeal_samples[41239]=5773;
squeal_samples[41240]=3544;
squeal_samples[41241]=5753;
squeal_samples[41242]=8577;
squeal_samples[41243]=11274;
squeal_samples[41244]=13856;
squeal_samples[41245]=16322;
squeal_samples[41246]=18674;
squeal_samples[41247]=20934;
squeal_samples[41248]=23082;
squeal_samples[41249]=25144;
squeal_samples[41250]=27108;
squeal_samples[41251]=28981;
squeal_samples[41252]=30785;
squeal_samples[41253]=32492;
squeal_samples[41254]=34135;
squeal_samples[41255]=35697;
squeal_samples[41256]=37187;
squeal_samples[41257]=38617;
squeal_samples[41258]=39976;
squeal_samples[41259]=41280;
squeal_samples[41260]=42521;
squeal_samples[41261]=43710;
squeal_samples[41262]=44839;
squeal_samples[41263]=45922;
squeal_samples[41264]=46957;
squeal_samples[41265]=47940;
squeal_samples[41266]=48884;
squeal_samples[41267]=49781;
squeal_samples[41268]=50642;
squeal_samples[41269]=51462;
squeal_samples[41270]=52249;
squeal_samples[41271]=52996;
squeal_samples[41272]=53713;
squeal_samples[41273]=54397;
squeal_samples[41274]=54569;
squeal_samples[41275]=49783;
squeal_samples[41276]=44006;
squeal_samples[41277]=38609;
squeal_samples[41278]=33545;
squeal_samples[41279]=28813;
squeal_samples[41280]=24379;
squeal_samples[41281]=20235;
squeal_samples[41282]=16353;
squeal_samples[41283]=12726;
squeal_samples[41284]=9319;
squeal_samples[41285]=6147;
squeal_samples[41286]=3577;
squeal_samples[41287]=5383;
squeal_samples[41288]=8226;
squeal_samples[41289]=10930;
squeal_samples[41290]=13533;
squeal_samples[41291]=16011;
squeal_samples[41292]=18373;
squeal_samples[41293]=20646;
squeal_samples[41294]=22807;
squeal_samples[41295]=24878;
squeal_samples[41296]=26858;
squeal_samples[41297]=28746;
squeal_samples[41298]=30554;
squeal_samples[41299]=32273;
squeal_samples[41300]=33924;
squeal_samples[41301]=35494;
squeal_samples[41302]=36998;
squeal_samples[41303]=38427;
squeal_samples[41304]=39803;
squeal_samples[41305]=41107;
squeal_samples[41306]=42364;
squeal_samples[41307]=43549;
squeal_samples[41308]=44697;
squeal_samples[41309]=45774;
squeal_samples[41310]=46821;
squeal_samples[41311]=47814;
squeal_samples[41312]=48755;
squeal_samples[41313]=49668;
squeal_samples[41314]=50523;
squeal_samples[41315]=51357;
squeal_samples[41316]=52139;
squeal_samples[41317]=52894;
squeal_samples[41318]=53615;
squeal_samples[41319]=54303;
squeal_samples[41320]=54914;
squeal_samples[41321]=51344;
squeal_samples[41322]=45478;
squeal_samples[41323]=39975;
squeal_samples[41324]=34834;
squeal_samples[41325]=30019;
squeal_samples[41326]=25503;
squeal_samples[41327]=21288;
squeal_samples[41328]=17340;
squeal_samples[41329]=13645;
squeal_samples[41330]=10188;
squeal_samples[41331]=6949;
squeal_samples[41332]=3963;
squeal_samples[41333]=4680;
squeal_samples[41334]=7543;
squeal_samples[41335]=10287;
squeal_samples[41336]=12914;
squeal_samples[41337]=15418;
squeal_samples[41338]=17813;
squeal_samples[41339]=20100;
squeal_samples[41340]=22294;
squeal_samples[41341]=24384;
squeal_samples[41342]=26386;
squeal_samples[41343]=28291;
squeal_samples[41344]=30123;
squeal_samples[41345]=31857;
squeal_samples[41346]=33532;
squeal_samples[41347]=35114;
squeal_samples[41348]=36638;
squeal_samples[41349]=38085;
squeal_samples[41350]=39469;
squeal_samples[41351]=40789;
squeal_samples[41352]=42061;
squeal_samples[41353]=43256;
squeal_samples[41354]=44421;
squeal_samples[41355]=45509;
squeal_samples[41356]=46569;
squeal_samples[41357]=47564;
squeal_samples[41358]=48531;
squeal_samples[41359]=49436;
squeal_samples[41360]=50322;
squeal_samples[41361]=51144;
squeal_samples[41362]=51948;
squeal_samples[41363]=52706;
squeal_samples[41364]=53440;
squeal_samples[41365]=54127;
squeal_samples[41366]=54799;
squeal_samples[41367]=52820;
squeal_samples[41368]=46904;
squeal_samples[41369]=41313;
squeal_samples[41370]=36086;
squeal_samples[41371]=31183;
squeal_samples[41372]=26606;
squeal_samples[41373]=22305;
squeal_samples[41374]=18298;
squeal_samples[41375]=14536;
squeal_samples[41376]=11025;
squeal_samples[41377]=7732;
squeal_samples[41378]=4650;
squeal_samples[41379]=3983;
squeal_samples[41380]=6832;
squeal_samples[41381]=9604;
squeal_samples[41382]=12261;
squeal_samples[41383]=14796;
squeal_samples[41384]=17221;
squeal_samples[41385]=19530;
squeal_samples[41386]=21748;
squeal_samples[41387]=23864;
squeal_samples[41388]=25880;
squeal_samples[41389]=27817;
squeal_samples[41390]=29657;
squeal_samples[41391]=31426;
squeal_samples[41392]=33108;
squeal_samples[41393]=34719;
squeal_samples[41394]=36249;
squeal_samples[41395]=37725;
squeal_samples[41396]=39120;
squeal_samples[41397]=40457;
squeal_samples[41398]=41738;
squeal_samples[41399]=42957;
squeal_samples[41400]=44124;
squeal_samples[41401]=45237;
squeal_samples[41402]=46300;
squeal_samples[41403]=47315;
squeal_samples[41404]=48282;
squeal_samples[41405]=49208;
squeal_samples[41406]=50090;
squeal_samples[41407]=50936;
squeal_samples[41408]=51741;
squeal_samples[41409]=52513;
squeal_samples[41410]=53247;
squeal_samples[41411]=53950;
squeal_samples[41412]=54628;
squeal_samples[41413]=53930;
squeal_samples[41414]=48351;
squeal_samples[41415]=42666;
squeal_samples[41416]=37350;
squeal_samples[41417]=32371;
squeal_samples[41418]=27709;
squeal_samples[41419]=23349;
squeal_samples[41420]=19260;
squeal_samples[41421]=15447;
squeal_samples[41422]=11872;
squeal_samples[41423]=8525;
squeal_samples[41424]=5392;
squeal_samples[41425]=3595;
squeal_samples[41426]=6111;
squeal_samples[41427]=8915;
squeal_samples[41428]=11598;
squeal_samples[41429]=14164;
squeal_samples[41430]=16610;
squeal_samples[41431]=18953;
squeal_samples[41432]=21194;
squeal_samples[41433]=23331;
squeal_samples[41434]=25380;
squeal_samples[41435]=27332;
squeal_samples[41436]=29198;
squeal_samples[41437]=30986;
squeal_samples[41438]=32681;
squeal_samples[41439]=34312;
squeal_samples[41440]=35865;
squeal_samples[41441]=37351;
squeal_samples[41442]=38762;
squeal_samples[41443]=40125;
squeal_samples[41444]=41408;
squeal_samples[41445]=42652;
squeal_samples[41446]=43825;
squeal_samples[41447]=44951;
squeal_samples[41448]=46023;
squeal_samples[41449]=47057;
squeal_samples[41450]=48029;
squeal_samples[41451]=48976;
squeal_samples[41452]=49857;
squeal_samples[41453]=50724;
squeal_samples[41454]=51532;
squeal_samples[41455]=52314;
squeal_samples[41456]=53056;
squeal_samples[41457]=53767;
squeal_samples[41458]=54447;
squeal_samples[41459]=54617;
squeal_samples[41460]=49822;
squeal_samples[41461]=44048;
squeal_samples[41462]=38637;
squeal_samples[41463]=33577;
squeal_samples[41464]=28836;
squeal_samples[41465]=24400;
squeal_samples[41466]=20246;
squeal_samples[41467]=16370;
squeal_samples[41468]=12730;
squeal_samples[41469]=9332;
squeal_samples[41470]=6146;
squeal_samples[41471]=3575;
squeal_samples[41472]=5383;
squeal_samples[41473]=8214;
squeal_samples[41474]=10927;
squeal_samples[41475]=13520;
squeal_samples[41476]=16002;
squeal_samples[41477]=18362;
squeal_samples[41478]=20634;
squeal_samples[41479]=22793;
squeal_samples[41480]=24865;
squeal_samples[41481]=26840;
squeal_samples[41482]=28726;
squeal_samples[41483]=30536;
squeal_samples[41484]=32253;
squeal_samples[41485]=33905;
squeal_samples[41486]=35473;
squeal_samples[41487]=36973;
squeal_samples[41488]=38411;
squeal_samples[41489]=39775;
squeal_samples[41490]=41091;
squeal_samples[41491]=42333;
squeal_samples[41492]=43531;
squeal_samples[41493]=44661;
squeal_samples[41494]=45756;
squeal_samples[41495]=46787;
squeal_samples[41496]=47786;
squeal_samples[41497]=48725;
squeal_samples[41498]=49638;
squeal_samples[41499]=50494;
squeal_samples[41500]=51328;
squeal_samples[41501]=52107;
squeal_samples[41502]=52866;
squeal_samples[41503]=53580;
squeal_samples[41504]=54273;
squeal_samples[41505]=54878;
squeal_samples[41506]=51317;
squeal_samples[41507]=45445;
squeal_samples[41508]=39948;
squeal_samples[41509]=34798;
squeal_samples[41510]=29982;
squeal_samples[41511]=25473;
squeal_samples[41512]=21248;
squeal_samples[41513]=17308;
squeal_samples[41514]=13602;
squeal_samples[41515]=10156;
squeal_samples[41516]=6911;
squeal_samples[41517]=3931;
squeal_samples[41518]=4642;
squeal_samples[41519]=7509;
squeal_samples[41520]=10254;
squeal_samples[41521]=12871;
squeal_samples[41522]=15379;
squeal_samples[41523]=17777;
squeal_samples[41524]=20065;
squeal_samples[41525]=22254;
squeal_samples[41526]=24350;
squeal_samples[41527]=26344;
squeal_samples[41528]=28258;
squeal_samples[41529]=30078;
squeal_samples[41530]=31823;
squeal_samples[41531]=33487;
squeal_samples[41532]=35076;
squeal_samples[41533]=36597;
squeal_samples[41534]=38043;
squeal_samples[41535]=39435;
squeal_samples[41536]=40752;
squeal_samples[41537]=42014;
squeal_samples[41538]=43228;
squeal_samples[41539]=44375;
squeal_samples[41540]=45478;
squeal_samples[41541]=46525;
squeal_samples[41542]=47528;
squeal_samples[41543]=48485;
squeal_samples[41544]=49402;
squeal_samples[41545]=50276;
squeal_samples[41546]=51106;
squeal_samples[41547]=51908;
squeal_samples[41548]=52665;
squeal_samples[41549]=53398;
squeal_samples[41550]=54095;
squeal_samples[41551]=54754;
squeal_samples[41552]=52784;
squeal_samples[41553]=46862;
squeal_samples[41554]=41278;
squeal_samples[41555]=36045;
squeal_samples[41556]=31143;
squeal_samples[41557]=26564;
squeal_samples[41558]=22269;
squeal_samples[41559]=18252;
squeal_samples[41560]=14501;
squeal_samples[41561]=10979;
squeal_samples[41562]=7698;
squeal_samples[41563]=4603;
squeal_samples[41564]=3948;
squeal_samples[41565]=6787;
squeal_samples[41566]=9567;
squeal_samples[41567]=12219;
squeal_samples[41568]=14757;
squeal_samples[41569]=17178;
squeal_samples[41570]=19492;
squeal_samples[41571]=21705;
squeal_samples[41572]=23825;
squeal_samples[41573]=25840;
squeal_samples[41574]=27776;
squeal_samples[41575]=29623;
squeal_samples[41576]=31383;
squeal_samples[41577]=33070;
squeal_samples[41578]=34676;
squeal_samples[41579]=36212;
squeal_samples[41580]=37681;
squeal_samples[41581]=39083;
squeal_samples[41582]=40420;
squeal_samples[41583]=41698;
squeal_samples[41584]=42916;
squeal_samples[41585]=44085;
squeal_samples[41586]=45196;
squeal_samples[41587]=46260;
squeal_samples[41588]=47274;
squeal_samples[41589]=48242;
squeal_samples[41590]=49167;
squeal_samples[41591]=50051;
squeal_samples[41592]=50895;
squeal_samples[41593]=51699;
squeal_samples[41594]=52475;
squeal_samples[41595]=53204;
squeal_samples[41596]=53912;
squeal_samples[41597]=54587;
squeal_samples[41598]=53889;
squeal_samples[41599]=48310;
squeal_samples[41600]=42627;
squeal_samples[41601]=37308;
squeal_samples[41602]=32332;
squeal_samples[41603]=27670;
squeal_samples[41604]=23305;
squeal_samples[41605]=19222;
squeal_samples[41606]=15406;
squeal_samples[41607]=11831;
squeal_samples[41608]=8487;
squeal_samples[41609]=5350;
squeal_samples[41610]=3554;
squeal_samples[41611]=6072;
squeal_samples[41612]=8873;
squeal_samples[41613]=11559;
squeal_samples[41614]=14123;
squeal_samples[41615]=16568;
squeal_samples[41616]=18916;
squeal_samples[41617]=21149;
squeal_samples[41618]=23295;
squeal_samples[41619]=25336;
squeal_samples[41620]=27293;
squeal_samples[41621]=29158;
squeal_samples[41622]=30945;
squeal_samples[41623]=32640;
squeal_samples[41624]=34271;
squeal_samples[41625]=35827;
squeal_samples[41626]=37308;
squeal_samples[41627]=38724;
squeal_samples[41628]=40081;
squeal_samples[41629]=41371;
squeal_samples[41630]=42609;
squeal_samples[41631]=43786;
squeal_samples[41632]=44908;
squeal_samples[41633]=45986;
squeal_samples[41634]=47013;
squeal_samples[41635]=47993;
squeal_samples[41636]=48929;
squeal_samples[41637]=49822;
squeal_samples[41638]=50679;
squeal_samples[41639]=51495;
squeal_samples[41640]=52271;
squeal_samples[41641]=53017;
squeal_samples[41642]=53724;
squeal_samples[41643]=54408;
squeal_samples[41644]=54846;
squeal_samples[41645]=50602;
squeal_samples[41646]=44780;
squeal_samples[41647]=39318;
squeal_samples[41648]=34211;
squeal_samples[41649]=29424;
squeal_samples[41650]=24952;
squeal_samples[41651]=20758;
squeal_samples[41652]=16846;
squeal_samples[41653]=13179;
squeal_samples[41654]=9741;
squeal_samples[41655]=6531;
squeal_samples[41656]=3707;
squeal_samples[41657]=5011;
squeal_samples[41658]=7858;
squeal_samples[41659]=10587;
squeal_samples[41660]=13194;
squeal_samples[41661]=15687;
squeal_samples[41662]=18058;
squeal_samples[41663]=20342;
squeal_samples[41664]=22514;
squeal_samples[41665]=24598;
squeal_samples[41666]=26579;
squeal_samples[41667]=28483;
squeal_samples[41668]=30291;
squeal_samples[41669]=32027;
squeal_samples[41670]=33677;
squeal_samples[41671]=35260;
squeal_samples[41672]=36764;
squeal_samples[41673]=38212;
squeal_samples[41674]=39585;
squeal_samples[41675]=40903;
squeal_samples[41676]=42152;
squeal_samples[41677]=43353;
squeal_samples[41678]=44498;
squeal_samples[41679]=45593;
squeal_samples[41680]=46636;
squeal_samples[41681]=47635;
squeal_samples[41682]=48582;
squeal_samples[41683]=49493;
squeal_samples[41684]=50357;
squeal_samples[41685]=51194;
squeal_samples[41686]=51981;
squeal_samples[41687]=52743;
squeal_samples[41688]=53461;
squeal_samples[41689]=54159;
squeal_samples[41690]=54816;
squeal_samples[41691]=52839;
squeal_samples[41692]=46914;
squeal_samples[41693]=41318;
squeal_samples[41694]=36086;
squeal_samples[41695]=31176;
squeal_samples[41696]=26596;
squeal_samples[41697]=22294;
squeal_samples[41698]=18275;
squeal_samples[41699]=14522;
squeal_samples[41700]=10994;
squeal_samples[41701]=7709;
squeal_samples[41702]=4619;
squeal_samples[41703]=3953;
squeal_samples[41704]=6796;
squeal_samples[41705]=9574;
squeal_samples[41706]=12221;
squeal_samples[41707]=14754;
squeal_samples[41708]=17181;
squeal_samples[41709]=19487;
squeal_samples[41710]=21704;
squeal_samples[41711]=23820;
squeal_samples[41712]=25838;
squeal_samples[41713]=27772;
squeal_samples[41714]=29614;
squeal_samples[41715]=31376;
squeal_samples[41716]=33060;
squeal_samples[41717]=34669;
squeal_samples[41718]=36200;
squeal_samples[41719]=37672;
squeal_samples[41720]=39062;
squeal_samples[41721]=40414;
squeal_samples[41722]=41676;
squeal_samples[41723]=42908;
squeal_samples[41724]=44062;
squeal_samples[41725]=45177;
squeal_samples[41726]=46241;
squeal_samples[41727]=47253;
squeal_samples[41728]=48223;
squeal_samples[41729]=49149;
squeal_samples[41730]=50029;
squeal_samples[41731]=50876;
squeal_samples[41732]=51680;
squeal_samples[41733]=52453;
squeal_samples[41734]=53188;
squeal_samples[41735]=53888;
squeal_samples[41736]=54563;
squeal_samples[41737]=54348;
squeal_samples[41738]=49100;
squeal_samples[41739]=43362;
squeal_samples[41740]=37995;
squeal_samples[41741]=32974;
squeal_samples[41742]=28264;
squeal_samples[41743]=23863;
squeal_samples[41744]=19738;
squeal_samples[41745]=15892;
squeal_samples[41746]=12279;
squeal_samples[41747]=8906;
squeal_samples[41748]=5745;
squeal_samples[41749]=3512;
squeal_samples[41750]=5720;
squeal_samples[41751]=8533;
squeal_samples[41752]=11231;
squeal_samples[41753]=13807;
squeal_samples[41754]=16277;
squeal_samples[41755]=18624;
squeal_samples[41756]=20874;
squeal_samples[41757]=23029;
squeal_samples[41758]=25082;
squeal_samples[41759]=27049;
squeal_samples[41760]=28918;
squeal_samples[41761]=30716;
squeal_samples[41762]=32426;
squeal_samples[41763]=34060;
squeal_samples[41764]=35624;
squeal_samples[41765]=37115;
squeal_samples[41766]=38541;
squeal_samples[41767]=39905;
squeal_samples[41768]=41200;
squeal_samples[41769]=42443;
squeal_samples[41770]=43626;
squeal_samples[41771]=44759;
squeal_samples[41772]=45838;
squeal_samples[41773]=46873;
squeal_samples[41774]=47851;
squeal_samples[41775]=48799;
squeal_samples[41776]=49691;
squeal_samples[41777]=50553;
squeal_samples[41778]=51369;
squeal_samples[41779]=52157;
squeal_samples[41780]=52903;
squeal_samples[41781]=53619;
squeal_samples[41782]=54306;
squeal_samples[41783]=54900;
squeal_samples[41784]=51342;
squeal_samples[41785]=45458;
squeal_samples[41786]=39958;
squeal_samples[41787]=34810;
squeal_samples[41788]=29984;
squeal_samples[41789]=25473;
squeal_samples[41790]=21242;
squeal_samples[41791]=17299;
squeal_samples[41792]=13595;
squeal_samples[41793]=10133;
squeal_samples[41794]=6899;
squeal_samples[41795]=3904;
squeal_samples[41796]=4623;
squeal_samples[41797]=7483;
squeal_samples[41798]=10229;
squeal_samples[41799]=12840;
squeal_samples[41800]=15354;
squeal_samples[41801]=17741;
squeal_samples[41802]=20033;
squeal_samples[41803]=22221;
squeal_samples[41804]=24309;
squeal_samples[41805]=26313;
squeal_samples[41806]=28218;
squeal_samples[41807]=30039;
squeal_samples[41808]=31785;
squeal_samples[41809]=33446;
squeal_samples[41810]=35040;
squeal_samples[41811]=36555;
squeal_samples[41812]=38008;
squeal_samples[41813]=39387;
squeal_samples[41814]=40715;
squeal_samples[41815]=41970;
squeal_samples[41816]=43176;
squeal_samples[41817]=44333;
squeal_samples[41818]=45427;
squeal_samples[41819]=46481;
squeal_samples[41820]=47479;
squeal_samples[41821]=48440;
squeal_samples[41822]=49351;
squeal_samples[41823]=50227;
squeal_samples[41824]=51057;
squeal_samples[41825]=51856;
squeal_samples[41826]=52618;
squeal_samples[41827]=53346;
squeal_samples[41828]=54038;
squeal_samples[41829]=54708;
squeal_samples[41830]=53413;
squeal_samples[41831]=47616;
squeal_samples[41832]=41963;
squeal_samples[41833]=36694;
squeal_samples[41834]=31742;
squeal_samples[41835]=27124;
squeal_samples[41836]=22787;
squeal_samples[41837]=18732;
squeal_samples[41838]=14948;
squeal_samples[41839]=11395;
squeal_samples[41840]=8076;
squeal_samples[41841]=4969;
squeal_samples[41842]=3684;
squeal_samples[41843]=6417;
squeal_samples[41844]=9198;
squeal_samples[41845]=11867;
squeal_samples[41846]=14413;
squeal_samples[41847]=16852;
squeal_samples[41848]=19176;
squeal_samples[41849]=21401;
squeal_samples[41850]=23530;
squeal_samples[41851]=25564;
squeal_samples[41852]=27502;
squeal_samples[41853]=29357;
squeal_samples[41854]=31133;
squeal_samples[41855]=32826;
squeal_samples[41856]=34440;
squeal_samples[41857]=35986;
squeal_samples[41858]=37455;
squeal_samples[41859]=38871;
squeal_samples[41860]=40209;
squeal_samples[41861]=41494;
squeal_samples[41862]=42723;
squeal_samples[41863]=43893;
squeal_samples[41864]=45008;
squeal_samples[41865]=46085;
squeal_samples[41866]=47093;
squeal_samples[41867]=48085;
squeal_samples[41868]=48998;
squeal_samples[41869]=49896;
squeal_samples[41870]=50739;
squeal_samples[41871]=51556;
squeal_samples[41872]=52322;
squeal_samples[41873]=53066;
squeal_samples[41874]=53771;
squeal_samples[41875]=54450;
squeal_samples[41876]=54612;
squeal_samples[41877]=49814;
squeal_samples[41878]=44032;
squeal_samples[41879]=38619;
squeal_samples[41880]=33548;
squeal_samples[41881]=28813;
squeal_samples[41882]=24367;
squeal_samples[41883]=20216;
squeal_samples[41884]=16328;
squeal_samples[41885]=12688;
squeal_samples[41886]=9285;
squeal_samples[41887]=6098;
squeal_samples[41888]=3529;
squeal_samples[41889]=5329;
squeal_samples[41890]=8161;
squeal_samples[41891]=10876;
squeal_samples[41892]=13460;
squeal_samples[41893]=15945;
squeal_samples[41894]=18298;
squeal_samples[41895]=20576;
squeal_samples[41896]=22729;
squeal_samples[41897]=24802;
squeal_samples[41898]=26774;
squeal_samples[41899]=28665;
squeal_samples[41900]=30465;
squeal_samples[41901]=32187;
squeal_samples[41902]=33827;
squeal_samples[41903]=35406;
squeal_samples[41904]=36904;
squeal_samples[41905]=38340;
squeal_samples[41906]=39704;
squeal_samples[41907]=41014;
squeal_samples[41908]=42261;
squeal_samples[41909]=43447;
squeal_samples[41910]=44592;
squeal_samples[41911]=45671;
squeal_samples[41912]=46716;
squeal_samples[41913]=47705;
squeal_samples[41914]=48650;
squeal_samples[41915]=49558;
squeal_samples[41916]=50416;
squeal_samples[41917]=51244;
squeal_samples[41918]=52032;
squeal_samples[41919]=52782;
squeal_samples[41920]=53501;
squeal_samples[41921]=54189;
squeal_samples[41922]=54849;
squeal_samples[41923]=52070;
squeal_samples[41924]=46148;
squeal_samples[41925]=40593;
squeal_samples[41926]=35406;
squeal_samples[41927]=30536;
squeal_samples[41928]=25989;
squeal_samples[41929]=21730;
squeal_samples[41930]=17741;
squeal_samples[41931]=14014;
squeal_samples[41932]=10523;
squeal_samples[41933]=7260;
squeal_samples[41934]=4200;
squeal_samples[41935]=4223;
squeal_samples[41936]=7100;
squeal_samples[41937]=9861;
squeal_samples[41938]=12491;
squeal_samples[41939]=15014;
squeal_samples[41940]=17422;
squeal_samples[41941]=19722;
squeal_samples[41942]=21924;
squeal_samples[41943]=24025;
squeal_samples[41944]=26037;
squeal_samples[41945]=27955;
squeal_samples[41946]=29787;
squeal_samples[41947]=31543;
squeal_samples[41948]=33210;
squeal_samples[41949]=34814;
squeal_samples[41950]=36336;
squeal_samples[41951]=37798;
squeal_samples[41952]=39189;
squeal_samples[41953]=40522;
squeal_samples[41954]=41788;
squeal_samples[41955]=43001;
squeal_samples[41956]=44160;
squeal_samples[41957]=45262;
squeal_samples[41958]=46321;
squeal_samples[41959]=47328;
squeal_samples[41960]=48292;
squeal_samples[41961]=49206;
squeal_samples[41962]=50089;
squeal_samples[41963]=50928;
squeal_samples[41964]=51729;
squeal_samples[41965]=52493;
squeal_samples[41966]=53225;
squeal_samples[41967]=53926;
squeal_samples[41968]=54592;
squeal_samples[41969]=54376;
squeal_samples[41970]=49118;
squeal_samples[41971]=43383;
squeal_samples[41972]=38012;
squeal_samples[41973]=32980;
squeal_samples[41974]=28277;
squeal_samples[41975]=23863;
squeal_samples[41976]=19741;
squeal_samples[41977]=15882;
squeal_samples[41978]=12274;
squeal_samples[41979]=8893;
squeal_samples[41980]=5732;
squeal_samples[41981]=3497;
squeal_samples[41982]=5700;
squeal_samples[41983]=8518;
squeal_samples[41984]=11210;
squeal_samples[41985]=13787;
squeal_samples[41986]=16252;
squeal_samples[41987]=18602;
squeal_samples[41988]=20851;
squeal_samples[41989]=23000;
squeal_samples[41990]=25055;
squeal_samples[41991]=27024;
squeal_samples[41992]=28892;
squeal_samples[41993]=30685;
squeal_samples[41994]=32398;
squeal_samples[41995]=34033;
squeal_samples[41996]=35594;
squeal_samples[41997]=37083;
squeal_samples[41998]=38506;
squeal_samples[41999]=39866;
squeal_samples[42000]=41164;
squeal_samples[42001]=42408;
squeal_samples[42002]=43587;
squeal_samples[42003]=44725;
squeal_samples[42004]=45795;
squeal_samples[42005]=46835;
squeal_samples[42006]=47811;
squeal_samples[42007]=48759;
squeal_samples[42008]=49655;
squeal_samples[42009]=50509;
squeal_samples[42010]=51335;
squeal_samples[42011]=52112;
squeal_samples[42012]=52862;
squeal_samples[42013]=53578;
squeal_samples[42014]=54259;
squeal_samples[42015]=54919;
squeal_samples[42016]=52134;
squeal_samples[42017]=46206;
squeal_samples[42018]=40642;
squeal_samples[42019]=35451;
squeal_samples[42020]=30583;
squeal_samples[42021]=26026;
squeal_samples[42022]=21767;
squeal_samples[42023]=17772;
squeal_samples[42024]=14045;
squeal_samples[42025]=10552;
squeal_samples[42026]=7281;
squeal_samples[42027]=4221;
squeal_samples[42028]=4238;
squeal_samples[42029]=7120;
squeal_samples[42030]=9872;
squeal_samples[42031]=12504;
squeal_samples[42032]=15026;
squeal_samples[42033]=17430;
squeal_samples[42034]=19734;
squeal_samples[42035]=21931;
squeal_samples[42036]=24031;
squeal_samples[42037]=26042;
squeal_samples[42038]=27959;
squeal_samples[42039]=29791;
squeal_samples[42040]=31543;
squeal_samples[42041]=33212;
squeal_samples[42042]=34816;
squeal_samples[42043]=36339;
squeal_samples[42044]=37791;
squeal_samples[42045]=39189;
squeal_samples[42046]=40515;
squeal_samples[42047]=41787;
squeal_samples[42048]=42995;
squeal_samples[42049]=44152;
squeal_samples[42050]=45258;
squeal_samples[42051]=46311;
squeal_samples[42052]=47321;
squeal_samples[42053]=48281;
squeal_samples[42054]=49203;
squeal_samples[42055]=50081;
squeal_samples[42056]=50916;
squeal_samples[42057]=51724;
squeal_samples[42058]=52481;
squeal_samples[42059]=53217;
squeal_samples[42060]=53912;
squeal_samples[42061]=54582;
squeal_samples[42062]=54363;
squeal_samples[42063]=49107;
squeal_samples[42064]=43371;
squeal_samples[42065]=37994;
squeal_samples[42066]=32969;
squeal_samples[42067]=28260;
squeal_samples[42068]=23850;
squeal_samples[42069]=19725;
squeal_samples[42070]=15870;
squeal_samples[42071]=12257;
squeal_samples[42072]=8881;
squeal_samples[42073]=5715;
squeal_samples[42074]=3485;
squeal_samples[42075]=5684;
squeal_samples[42076]=8504;
squeal_samples[42077]=11196;
squeal_samples[42078]=13772;
squeal_samples[42079]=16233;
squeal_samples[42080]=18581;
squeal_samples[42081]=20837;
squeal_samples[42082]=22984;
squeal_samples[42083]=25039;
squeal_samples[42084]=26999;
squeal_samples[42085]=28882;
squeal_samples[42086]=30666;
squeal_samples[42087]=32383;
squeal_samples[42088]=34009;
squeal_samples[42089]=35576;
squeal_samples[42090]=37068;
squeal_samples[42091]=38485;
squeal_samples[42092]=39855;
squeal_samples[42093]=41141;
squeal_samples[42094]=42394;
squeal_samples[42095]=43568;
squeal_samples[42096]=44703;
squeal_samples[42097]=45779;
squeal_samples[42098]=46813;
squeal_samples[42099]=47797;
squeal_samples[42100]=48739;
squeal_samples[42101]=49633;
squeal_samples[42102]=50493;
squeal_samples[42103]=51311;
squeal_samples[42104]=52097;
squeal_samples[42105]=52842;
squeal_samples[42106]=53563;
squeal_samples[42107]=54236;
squeal_samples[42108]=54901;
squeal_samples[42109]=52113;
squeal_samples[42110]=46186;
squeal_samples[42111]=40629;
squeal_samples[42112]=35431;
squeal_samples[42113]=30561;
squeal_samples[42114]=26010;
squeal_samples[42115]=21743;
squeal_samples[42116]=17755;
squeal_samples[42117]=14025;
squeal_samples[42118]=10530;
squeal_samples[42119]=7264;
squeal_samples[42120]=4199;
squeal_samples[42121]=4220;
squeal_samples[42122]=7099;
squeal_samples[42123]=9858;
squeal_samples[42124]=12484;
squeal_samples[42125]=15007;
squeal_samples[42126]=17409;
squeal_samples[42127]=19715;
squeal_samples[42128]=21910;
squeal_samples[42129]=24014;
squeal_samples[42130]=26019;
squeal_samples[42131]=27941;
squeal_samples[42132]=29771;
squeal_samples[42133]=31521;
squeal_samples[42134]=33196;
squeal_samples[42135]=34793;
squeal_samples[42136]=36320;
squeal_samples[42137]=37773;
squeal_samples[42138]=39166;
squeal_samples[42139]=40499;
squeal_samples[42140]=41762;
squeal_samples[42141]=42980;
squeal_samples[42142]=44129;
squeal_samples[42143]=45240;
squeal_samples[42144]=46291;
squeal_samples[42145]=47300;
squeal_samples[42146]=48262;
squeal_samples[42147]=49183;
squeal_samples[42148]=50061;
squeal_samples[42149]=50897;
squeal_samples[42150]=51703;
squeal_samples[42151]=52462;
squeal_samples[42152]=53197;
squeal_samples[42153]=53891;
squeal_samples[42154]=54564;
squeal_samples[42155]=54341;
squeal_samples[42156]=49090;
squeal_samples[42157]=43348;
squeal_samples[42158]=37977;
squeal_samples[42159]=32947;
squeal_samples[42160]=28241;
squeal_samples[42161]=23831;
squeal_samples[42162]=19704;
squeal_samples[42163]=15851;
squeal_samples[42164]=12236;
squeal_samples[42165]=8861;
squeal_samples[42166]=5699;
squeal_samples[42167]=3460;
squeal_samples[42168]=5669;
squeal_samples[42169]=8480;
squeal_samples[42170]=11178;
squeal_samples[42171]=13754;
squeal_samples[42172]=16209;
squeal_samples[42173]=18567;
squeal_samples[42174]=20812;
squeal_samples[42175]=22969;
squeal_samples[42176]=25014;
squeal_samples[42177]=26984;
squeal_samples[42178]=28859;
squeal_samples[42179]=30650;
squeal_samples[42180]=32359;
squeal_samples[42181]=33993;
squeal_samples[42182]=35554;
squeal_samples[42183]=37049;
squeal_samples[42184]=38467;
squeal_samples[42185]=39830;
squeal_samples[42186]=41128;
squeal_samples[42187]=42368;
squeal_samples[42188]=43553;
squeal_samples[42189]=44680;
squeal_samples[42190]=45762;
squeal_samples[42191]=46789;
squeal_samples[42192]=47781;
squeal_samples[42193]=48718;
squeal_samples[42194]=49613;
squeal_samples[42195]=50475;
squeal_samples[42196]=51289;
squeal_samples[42197]=52079;
squeal_samples[42198]=52821;
squeal_samples[42199]=53544;
squeal_samples[42200]=54217;
squeal_samples[42201]=54879;
squeal_samples[42202]=52097;
squeal_samples[42203]=46162;
squeal_samples[42204]=40612;
squeal_samples[42205]=35410;
squeal_samples[42206]=30542;
squeal_samples[42207]=25989;
squeal_samples[42208]=21725;
squeal_samples[42209]=17734;
squeal_samples[42210]=14005;
squeal_samples[42211]=10512;
squeal_samples[42212]=7242;
squeal_samples[42213]=4181;
squeal_samples[42214]=4199;
squeal_samples[42215]=7081;
squeal_samples[42216]=9836;
squeal_samples[42217]=12467;
squeal_samples[42218]=14984;
squeal_samples[42219]=17393;
squeal_samples[42220]=19693;
squeal_samples[42221]=21891;
squeal_samples[42222]=23993;
squeal_samples[42223]=26001;
squeal_samples[42224]=27921;
squeal_samples[42225]=29750;
squeal_samples[42226]=31504;
squeal_samples[42227]=33172;
squeal_samples[42228]=34778;
squeal_samples[42229]=36297;
squeal_samples[42230]=37754;
squeal_samples[42231]=39147;
squeal_samples[42232]=40477;
squeal_samples[42233]=41747;
squeal_samples[42234]=42956;
squeal_samples[42235]=44112;
squeal_samples[42236]=45218;
squeal_samples[42237]=46273;
squeal_samples[42238]=47279;
squeal_samples[42239]=48243;
squeal_samples[42240]=49164;
squeal_samples[42241]=50040;
squeal_samples[42242]=50879;
squeal_samples[42243]=51682;
squeal_samples[42244]=52442;
squeal_samples[42245]=53179;
squeal_samples[42246]=53870;
squeal_samples[42247]=54546;
squeal_samples[42248]=54319;
squeal_samples[42249]=49072;
squeal_samples[42250]=43329;
squeal_samples[42251]=37955;
squeal_samples[42252]=32930;
squeal_samples[42253]=28219;
squeal_samples[42254]=23812;
squeal_samples[42255]=19686;
squeal_samples[42256]=15828;
squeal_samples[42257]=12220;
squeal_samples[42258]=8839;
squeal_samples[42259]=5679;
squeal_samples[42260]=3442;
squeal_samples[42261]=5647;
squeal_samples[42262]=8463;
squeal_samples[42263]=11156;
squeal_samples[42264]=13735;
squeal_samples[42265]=16190;
squeal_samples[42266]=18545;
squeal_samples[42267]=20796;
squeal_samples[42268]=22945;
squeal_samples[42269]=24999;
squeal_samples[42270]=26960;
squeal_samples[42271]=28842;
squeal_samples[42272]=30628;
squeal_samples[42273]=32342;
squeal_samples[42274]=33971;
squeal_samples[42275]=35536;
squeal_samples[42276]=37028;
squeal_samples[42277]=38447;
squeal_samples[42278]=39813;
squeal_samples[42279]=41105;
squeal_samples[42280]=42351;
squeal_samples[42281]=43532;
squeal_samples[42282]=44661;
squeal_samples[42283]=45740;
squeal_samples[42284]=46773;
squeal_samples[42285]=47759;
squeal_samples[42286]=48699;
squeal_samples[42287]=49594;
squeal_samples[42288]=50452;
squeal_samples[42289]=51274;
squeal_samples[42290]=52054;
squeal_samples[42291]=52809;
squeal_samples[42292]=53515;
squeal_samples[42293]=54205;
squeal_samples[42294]=54855;
squeal_samples[42295]=52078;
squeal_samples[42296]=46144;
squeal_samples[42297]=40592;
squeal_samples[42298]=35389;
squeal_samples[42299]=30525;
squeal_samples[42300]=25966;
squeal_samples[42301]=21706;
squeal_samples[42302]=17717;
squeal_samples[42303]=13983;
squeal_samples[42304]=10494;
squeal_samples[42305]=7221;
squeal_samples[42306]=4161;
squeal_samples[42307]=4181;
squeal_samples[42308]=7059;
squeal_samples[42309]=9819;
squeal_samples[42310]=12444;
squeal_samples[42311]=14968;
squeal_samples[42312]=17370;
squeal_samples[42313]=19676;
squeal_samples[42314]=21869;
squeal_samples[42315]=23976;
squeal_samples[42316]=25977;
squeal_samples[42317]=27906;
squeal_samples[42318]=29727;
squeal_samples[42319]=31487;
squeal_samples[42320]=33151;
squeal_samples[42321]=34758;
squeal_samples[42322]=36277;
squeal_samples[42323]=37736;
squeal_samples[42324]=39126;
squeal_samples[42325]=40459;
squeal_samples[42326]=41725;
squeal_samples[42327]=42938;
squeal_samples[42328]=44091;
squeal_samples[42329]=45200;
squeal_samples[42330]=46251;
squeal_samples[42331]=47262;
squeal_samples[42332]=48221;
squeal_samples[42333]=49145;
squeal_samples[42334]=50020;
squeal_samples[42335]=50859;
squeal_samples[42336]=51661;
squeal_samples[42337]=52425;
squeal_samples[42338]=53156;
squeal_samples[42339]=53851;
squeal_samples[42340]=54525;
squeal_samples[42341]=54675;
squeal_samples[42342]=49866;
squeal_samples[42343]=44075;
squeal_samples[42344]=38654;
squeal_samples[42345]=33576;
squeal_samples[42346]=28825;
squeal_samples[42347]=24379;
squeal_samples[42348]=20217;
squeal_samples[42349]=16329;
squeal_samples[42350]=12679;
squeal_samples[42351]=9274;
squeal_samples[42352]=6074;
squeal_samples[42353]=3501;
squeal_samples[42354]=5299;
squeal_samples[42355]=8129;
squeal_samples[42356]=10838;
squeal_samples[42357]=13426;
squeal_samples[42358]=15900;
squeal_samples[42359]=18264;
squeal_samples[42360]=20526;
squeal_samples[42361]=22689;
squeal_samples[42362]=24747;
squeal_samples[42363]=26728;
squeal_samples[42364]=28606;
squeal_samples[42365]=30412;
squeal_samples[42366]=32129;
squeal_samples[42367]=33774;
squeal_samples[42368]=35342;
squeal_samples[42369]=36840;
squeal_samples[42370]=38271;
squeal_samples[42371]=39640;
squeal_samples[42372]=40939;
squeal_samples[42373]=42191;
squeal_samples[42374]=43381;
squeal_samples[42375]=44518;
squeal_samples[42376]=45601;
squeal_samples[42377]=46636;
squeal_samples[42378]=47635;
squeal_samples[42379]=48571;
squeal_samples[42380]=49482;
squeal_samples[42381]=50337;
squeal_samples[42382]=51162;
squeal_samples[42383]=51949;
squeal_samples[42384]=52697;
squeal_samples[42385]=53419;
squeal_samples[42386]=54104;
squeal_samples[42387]=54760;
squeal_samples[42388]=53466;
squeal_samples[42389]=47645;
squeal_samples[42390]=41994;
squeal_samples[42391]=36707;
squeal_samples[42392]=31750;
squeal_samples[42393]=27124;
squeal_samples[42394]=22782;
squeal_samples[42395]=18722;
squeal_samples[42396]=14926;
squeal_samples[42397]=11367;
squeal_samples[42398]=8041;
squeal_samples[42399]=4930;
squeal_samples[42400]=3643;
squeal_samples[42401]=6366;
squeal_samples[42402]=9151;
squeal_samples[42403]=11813;
squeal_samples[42404]=14359;
squeal_samples[42405]=16794;
squeal_samples[42406]=19115;
squeal_samples[42407]=21338;
squeal_samples[42408]=23464;
squeal_samples[42409]=25494;
squeal_samples[42410]=27433;
squeal_samples[42411]=29286;
squeal_samples[42412]=31059;
squeal_samples[42413]=32741;
squeal_samples[42414]=34364;
squeal_samples[42415]=35900;
squeal_samples[42416]=37379;
squeal_samples[42417]=38782;
squeal_samples[42418]=40128;
squeal_samples[42419]=41409;
squeal_samples[42420]=42634;
squeal_samples[42421]=43808;
squeal_samples[42422]=44918;
squeal_samples[42423]=45989;
squeal_samples[42424]=47006;
squeal_samples[42425]=47983;
squeal_samples[42426]=48904;
squeal_samples[42427]=49802;
squeal_samples[42428]=50644;
squeal_samples[42429]=51455;
squeal_samples[42430]=52227;
squeal_samples[42431]=52967;
squeal_samples[42432]=53669;
squeal_samples[42433]=54346;
squeal_samples[42434]=54938;
squeal_samples[42435]=51361;
squeal_samples[42436]=45474;
squeal_samples[42437]=39966;
squeal_samples[42438]=34798;
squeal_samples[42439]=29975;
squeal_samples[42440]=25448;
squeal_samples[42441]=21216;
squeal_samples[42442]=17263;
squeal_samples[42443]=13551;
squeal_samples[42444]=10090;
squeal_samples[42445]=6837;
squeal_samples[42446]=3852;
squeal_samples[42447]=4556;
squeal_samples[42448]=7418;
squeal_samples[42449]=10157;
squeal_samples[42450]=12775;
squeal_samples[42451]=15279;
squeal_samples[42452]=17662;
squeal_samples[42453]=19954;
squeal_samples[42454]=22135;
squeal_samples[42455]=24227;
squeal_samples[42456]=26222;
squeal_samples[42457]=28127;
squeal_samples[42458]=29952;
squeal_samples[42459]=31686;
squeal_samples[42460]=33354;
squeal_samples[42461]=34936;
squeal_samples[42462]=36458;
squeal_samples[42463]=37898;
squeal_samples[42464]=39284;
squeal_samples[42465]=40607;
squeal_samples[42466]=41864;
squeal_samples[42467]=43071;
squeal_samples[42468]=44220;
squeal_samples[42469]=45316;
squeal_samples[42470]=46364;
squeal_samples[42471]=47367;
squeal_samples[42472]=48322;
squeal_samples[42473]=49236;
squeal_samples[42474]=50108;
squeal_samples[42475]=50940;
squeal_samples[42476]=51740;
squeal_samples[42477]=52498;
squeal_samples[42478]=53225;
squeal_samples[42479]=53914;
squeal_samples[42480]=54584;
squeal_samples[42481]=54355;
squeal_samples[42482]=49102;
squeal_samples[42483]=43352;
squeal_samples[42484]=37980;
squeal_samples[42485]=32944;
squeal_samples[42486]=28231;
squeal_samples[42487]=23821;
squeal_samples[42488]=19693;
squeal_samples[42489]=15831;
squeal_samples[42490]=12223;
squeal_samples[42491]=8830;
squeal_samples[42492]=5670;
squeal_samples[42493]=3430;
squeal_samples[42494]=5636;
squeal_samples[42495]=8446;
squeal_samples[42496]=11141;
squeal_samples[42497]=13717;
squeal_samples[42498]=16175;
squeal_samples[42499]=18528;
squeal_samples[42500]=20773;
squeal_samples[42501]=22924;
squeal_samples[42502]=24977;
squeal_samples[42503]=26939;
squeal_samples[42504]=28813;
squeal_samples[42505]=30603;
squeal_samples[42506]=32312;
squeal_samples[42507]=33946;
squeal_samples[42508]=35502;
squeal_samples[42509]=36995;
squeal_samples[42510]=38415;
squeal_samples[42511]=39780;
squeal_samples[42512]=41072;
squeal_samples[42513]=42314;
squeal_samples[42514]=43497;
squeal_samples[42515]=44630;
squeal_samples[42516]=45707;
squeal_samples[42517]=46740;
squeal_samples[42518]=47720;
squeal_samples[42519]=48662;
squeal_samples[42520]=49554;
squeal_samples[42521]=50417;
squeal_samples[42522]=51232;
squeal_samples[42523]=52019;
squeal_samples[42524]=52760;
squeal_samples[42525]=53478;
squeal_samples[42526]=54159;
squeal_samples[42527]=54816;
squeal_samples[42528]=52826;
squeal_samples[42529]=46893;
squeal_samples[42530]=41287;
squeal_samples[42531]=36040;
squeal_samples[42532]=31133;
squeal_samples[42533]=26531;
squeal_samples[42534]=22235;
squeal_samples[42535]=18200;
squeal_samples[42536]=14444;
squeal_samples[42537]=10907;
squeal_samples[42538]=7617;
squeal_samples[42539]=4522;
squeal_samples[42540]=3851;
squeal_samples[42541]=6688;
squeal_samples[42542]=9465;
squeal_samples[42543]=12110;
squeal_samples[42544]=14638;
squeal_samples[42545]=17064;
squeal_samples[42546]=19369;
squeal_samples[42547]=21578;
squeal_samples[42548]=23698;
squeal_samples[42549]=25713;
squeal_samples[42550]=27642;
squeal_samples[42551]=29481;
squeal_samples[42552]=31244;
squeal_samples[42553]=32922;
squeal_samples[42554]=34526;
squeal_samples[42555]=36064;
squeal_samples[42556]=37526;
squeal_samples[42557]=38928;
squeal_samples[42558]=40262;
squeal_samples[42559]=41535;
squeal_samples[42560]=42754;
squeal_samples[42561]=43917;
squeal_samples[42562]=45032;
squeal_samples[42563]=46088;
squeal_samples[42564]=47105;
squeal_samples[42565]=48068;
squeal_samples[42566]=48995;
squeal_samples[42567]=49870;
squeal_samples[42568]=50722;
squeal_samples[42569]=51521;
squeal_samples[42570]=52293;
squeal_samples[42571]=53022;
squeal_samples[42572]=53729;
squeal_samples[42573]=54397;
squeal_samples[42574]=54828;
squeal_samples[42575]=50579;
squeal_samples[42576]=44735;
squeal_samples[42577]=39271;
squeal_samples[42578]=34148;
squeal_samples[42579]=29367;
squeal_samples[42580]=24875;
squeal_samples[42581]=20681;
squeal_samples[42582]=16756;
squeal_samples[42583]=13076;
squeal_samples[42584]=9644;
squeal_samples[42585]=6416;
squeal_samples[42586]=3594;
squeal_samples[42587]=4891;
squeal_samples[42588]=7737;
squeal_samples[42589]=10458;
squeal_samples[42590]=13063;
squeal_samples[42591]=15551;
squeal_samples[42592]=17929;
squeal_samples[42593]=20199;
squeal_samples[42594]=22374;
squeal_samples[42595]=24451;
squeal_samples[42596]=26437;
squeal_samples[42597]=28332;
squeal_samples[42598]=30145;
squeal_samples[42599]=31868;
squeal_samples[42600]=33527;
squeal_samples[42601]=35100;
squeal_samples[42602]=36614;
squeal_samples[42603]=38048;
squeal_samples[42604]=39423;
squeal_samples[42605]=40734;
squeal_samples[42606]=41989;
squeal_samples[42607]=43186;
squeal_samples[42608]=44332;
squeal_samples[42609]=45424;
squeal_samples[42610]=46462;
squeal_samples[42611]=47461;
squeal_samples[42612]=48410;
squeal_samples[42613]=49320;
squeal_samples[42614]=50190;
squeal_samples[42615]=51011;
squeal_samples[42616]=51811;
squeal_samples[42617]=52560;
squeal_samples[42618]=53283;
squeal_samples[42619]=53974;
squeal_samples[42620]=54633;
squeal_samples[42621]=53930;
squeal_samples[42622]=48327;
squeal_samples[42623]=42638;
squeal_samples[42624]=37301;
squeal_samples[42625]=32308;
squeal_samples[42626]=27632;
squeal_samples[42627]=23260;
squeal_samples[42628]=19167;
squeal_samples[42629]=15339;
squeal_samples[42630]=11754;
squeal_samples[42631]=8399;
squeal_samples[42632]=5255;
squeal_samples[42633]=3453;
squeal_samples[42634]=5964;
squeal_samples[42635]=8767;
squeal_samples[42636]=11436;
squeal_samples[42637]=14003;
squeal_samples[42638]=16443;
squeal_samples[42639]=18782;
squeal_samples[42640]=21016;
squeal_samples[42641]=23155;
squeal_samples[42642]=25197;
squeal_samples[42643]=27147;
squeal_samples[42644]=29014;
squeal_samples[42645]=30789;
squeal_samples[42646]=32489;
squeal_samples[42647]=34119;
squeal_samples[42648]=35665;
squeal_samples[42649]=37153;
squeal_samples[42650]=38559;
squeal_samples[42651]=39910;
squeal_samples[42652]=41206;
squeal_samples[42653]=42430;
squeal_samples[42654]=43614;
squeal_samples[42655]=44733;
squeal_samples[42656]=45810;
squeal_samples[42657]=46834;
squeal_samples[42658]=47811;
squeal_samples[42659]=48746;
squeal_samples[42660]=49639;
squeal_samples[42661]=50495;
squeal_samples[42662]=51303;
squeal_samples[42663]=52079;
squeal_samples[42664]=52826;
squeal_samples[42665]=53532;
squeal_samples[42666]=54214;
squeal_samples[42667]=54866;
squeal_samples[42668]=52868;
squeal_samples[42669]=46936;
squeal_samples[42670]=41320;
squeal_samples[42671]=36073;
squeal_samples[42672]=31155;
squeal_samples[42673]=26558;
squeal_samples[42674]=22253;
squeal_samples[42675]=18222;
squeal_samples[42676]=14454;
squeal_samples[42677]=10926;
squeal_samples[42678]=7620;
squeal_samples[42679]=4532;
squeal_samples[42680]=3846;
squeal_samples[42681]=6699;
squeal_samples[42682]=9463;
squeal_samples[42683]=12115;
squeal_samples[42684]=14643;
squeal_samples[42685]=17059;
squeal_samples[42686]=19368;
squeal_samples[42687]=21576;
squeal_samples[42688]=23689;
squeal_samples[42689]=25706;
squeal_samples[42690]=27636;
squeal_samples[42691]=29469;
squeal_samples[42692]=31236;
squeal_samples[42693]=32909;
squeal_samples[42694]=34523;
squeal_samples[42695]=36047;
squeal_samples[42696]=37516;
squeal_samples[42697]=38913;
squeal_samples[42698]=40249;
squeal_samples[42699]=41523;
squeal_samples[42700]=42740;
squeal_samples[42701]=43899;
squeal_samples[42702]=45013;
squeal_samples[42703]=46069;
squeal_samples[42704]=47087;
squeal_samples[42705]=48050;
squeal_samples[42706]=48975;
squeal_samples[42707]=49853;
squeal_samples[42708]=50695;
squeal_samples[42709]=51500;
squeal_samples[42710]=52272;
squeal_samples[42711]=53004;
squeal_samples[42712]=53711;
squeal_samples[42713]=54375;
squeal_samples[42714]=54971;
squeal_samples[42715]=51380;
squeal_samples[42716]=45495;
squeal_samples[42717]=39973;
squeal_samples[42718]=34815;
squeal_samples[42719]=29972;
squeal_samples[42720]=25453;
squeal_samples[42721]=21208;
squeal_samples[42722]=17254;
squeal_samples[42723]=13542;
squeal_samples[42724]=10074;
squeal_samples[42725]=6824;
squeal_samples[42726]=3828;
squeal_samples[42727]=4532;
squeal_samples[42728]=7391;
squeal_samples[42729]=10132;
squeal_samples[42730]=12747;
squeal_samples[42731]=15250;
squeal_samples[42732]=17633;
squeal_samples[42733]=19926;
squeal_samples[42734]=22101;
squeal_samples[42735]=24197;
squeal_samples[42736]=26182;
squeal_samples[42737]=28100;
squeal_samples[42738]=29910;
squeal_samples[42739]=31653;
squeal_samples[42740]=33310;
squeal_samples[42741]=34900;
squeal_samples[42742]=36414;
squeal_samples[42743]=37863;
squeal_samples[42744]=39239;
squeal_samples[42745]=40567;
squeal_samples[42746]=41821;
squeal_samples[42747]=43029;
squeal_samples[42748]=44172;
squeal_samples[42749]=45273;
squeal_samples[42750]=46323;
squeal_samples[42751]=47318;
squeal_samples[42752]=48275;
squeal_samples[42753]=49188;
squeal_samples[42754]=50060;
squeal_samples[42755]=50893;
squeal_samples[42756]=51691;
squeal_samples[42757]=52445;
squeal_samples[42758]=53178;
squeal_samples[42759]=53864;
squeal_samples[42760]=54537;
squeal_samples[42761]=54677;
squeal_samples[42762]=49866;
squeal_samples[42763]=44069;
squeal_samples[42764]=38640;
squeal_samples[42765]=33567;
squeal_samples[42766]=28805;
squeal_samples[42767]=24357;
squeal_samples[42768]=20184;
squeal_samples[42769]=16294;
squeal_samples[42770]=12642;
squeal_samples[42771]=9233;
squeal_samples[42772]=6036;
squeal_samples[42773]=3455;
squeal_samples[42774]=5251;
squeal_samples[42775]=8077;
squeal_samples[42776]=10786;
squeal_samples[42777]=13371;
squeal_samples[42778]=15850;
squeal_samples[42779]=18203;
squeal_samples[42780]=20470;
squeal_samples[42781]=22625;
squeal_samples[42782]=24689;
squeal_samples[42783]=26665;
squeal_samples[42784]=28547;
squeal_samples[42785]=30343;
squeal_samples[42786]=32067;
squeal_samples[42787]=33703;
squeal_samples[42788]=35281;
squeal_samples[42789]=36768;
squeal_samples[42790]=38210;
squeal_samples[42791]=39565;
squeal_samples[42792]=40875;
squeal_samples[42793]=42117;
squeal_samples[42794]=43311;
squeal_samples[42795]=44444;
squeal_samples[42796]=45532;
squeal_samples[42797]=46564;
squeal_samples[42798]=47556;
squeal_samples[42799]=48497;
squeal_samples[42800]=49401;
squeal_samples[42801]=50262;
squeal_samples[42802]=51085;
squeal_samples[42803]=51870;
squeal_samples[42804]=52622;
squeal_samples[42805]=53340;
squeal_samples[42806]=54027;
squeal_samples[42807]=54683;
squeal_samples[42808]=53968;
squeal_samples[42809]=48373;
squeal_samples[42810]=42666;
squeal_samples[42811]=37330;
squeal_samples[42812]=32333;
squeal_samples[42813]=27657;
squeal_samples[42814]=23276;
squeal_samples[42815]=19177;
squeal_samples[42816]=15348;
squeal_samples[42817]=11758;
squeal_samples[42818]=8404;
squeal_samples[42819]=5259;
squeal_samples[42820]=3453;
squeal_samples[42821]=5956;
squeal_samples[42822]=8760;
squeal_samples[42823]=11430;
squeal_samples[42824]=13997;
squeal_samples[42825]=16436;
squeal_samples[42826]=18777;
squeal_samples[42827]=21000;
squeal_samples[42828]=23148;
squeal_samples[42829]=25180;
squeal_samples[42830]=27136;
squeal_samples[42831]=28990;
squeal_samples[42832]=30777;
squeal_samples[42833]=32468;
squeal_samples[42834]=34098;
squeal_samples[42835]=35642;
squeal_samples[42836]=37131;
squeal_samples[42837]=38539;
squeal_samples[42838]=39892;
squeal_samples[42839]=41177;
squeal_samples[42840]=42413;
squeal_samples[42841]=43588;
squeal_samples[42842]=44712;
squeal_samples[42843]=45780;
squeal_samples[42844]=46807;
squeal_samples[42845]=47783;
squeal_samples[42846]=48716;
squeal_samples[42847]=49614;
squeal_samples[42848]=50459;
squeal_samples[42849]=51275;
squeal_samples[42850]=52051;
squeal_samples[42851]=52798;
squeal_samples[42852]=53503;
squeal_samples[42853]=54183;
squeal_samples[42854]=54830;
squeal_samples[42855]=52841;
squeal_samples[42856]=46901;
squeal_samples[42857]=41288;
squeal_samples[42858]=36044;
squeal_samples[42859]=31122;
squeal_samples[42860]=26525;
squeal_samples[42861]=22218;
squeal_samples[42862]=18184;
squeal_samples[42863]=14421;
squeal_samples[42864]=10890;
squeal_samples[42865]=7590;
squeal_samples[42866]=4494;
squeal_samples[42867]=3817;
squeal_samples[42868]=6663;
squeal_samples[42869]=9424;
squeal_samples[42870]=12078;
squeal_samples[42871]=14600;
squeal_samples[42872]=17030;
squeal_samples[42873]=19326;
squeal_samples[42874]=21539;
squeal_samples[42875]=23649;
squeal_samples[42876]=25667;
squeal_samples[42877]=27597;
squeal_samples[42878]=29438;
squeal_samples[42879]=31198;
squeal_samples[42880]=32875;
squeal_samples[42881]=34479;
squeal_samples[42882]=36012;
squeal_samples[42883]=37475;
squeal_samples[42884]=38874;
squeal_samples[42885]=40210;
squeal_samples[42886]=41486;
squeal_samples[42887]=42697;
squeal_samples[42888]=43865;
squeal_samples[42889]=44969;
squeal_samples[42890]=46035;
squeal_samples[42891]=47044;
squeal_samples[42892]=48013;
squeal_samples[42893]=48936;
squeal_samples[42894]=49818;
squeal_samples[42895]=50664;
squeal_samples[42896]=51464;
squeal_samples[42897]=52234;
squeal_samples[42898]=52966;
squeal_samples[42899]=53670;
squeal_samples[42900]=54338;
squeal_samples[42901]=54929;
squeal_samples[42902]=51345;
squeal_samples[42903]=45452;
squeal_samples[42904]=39938;
squeal_samples[42905]=34772;
squeal_samples[42906]=29937;
squeal_samples[42907]=25410;
squeal_samples[42908]=21178;
squeal_samples[42909]=17213;
squeal_samples[42910]=13504;
squeal_samples[42911]=10034;
squeal_samples[42912]=6786;
squeal_samples[42913]=3788;
squeal_samples[42914]=4495;
squeal_samples[42915]=7350;
squeal_samples[42916]=10094;
squeal_samples[42917]=12709;
squeal_samples[42918]=15208;
squeal_samples[42919]=17599;
squeal_samples[42920]=19880;
squeal_samples[42921]=22070;
squeal_samples[42922]=24151;
squeal_samples[42923]=26149;
squeal_samples[42924]=28056;
squeal_samples[42925]=29874;
squeal_samples[42926]=31613;
squeal_samples[42927]=33277;
squeal_samples[42928]=34860;
squeal_samples[42929]=36376;
squeal_samples[42930]=37824;
squeal_samples[42931]=39199;
squeal_samples[42932]=40530;
squeal_samples[42933]=41779;
squeal_samples[42934]=42993;
squeal_samples[42935]=44136;
squeal_samples[42936]=45237;
squeal_samples[42937]=46280;
squeal_samples[42938]=47282;
squeal_samples[42939]=48235;
squeal_samples[42940]=49149;
squeal_samples[42941]=50022;
squeal_samples[42942]=50852;
squeal_samples[42943]=51653;
squeal_samples[42944]=52406;
squeal_samples[42945]=53138;
squeal_samples[42946]=53828;
squeal_samples[42947]=54495;
squeal_samples[42948]=54639;
squeal_samples[42949]=49829;
squeal_samples[42950]=44025;
squeal_samples[42951]=38607;
squeal_samples[42952]=33522;
squeal_samples[42953]=28772;
squeal_samples[42954]=24314;
squeal_samples[42955]=20147;
squeal_samples[42956]=16254;
squeal_samples[42957]=12602;
squeal_samples[42958]=9195;
squeal_samples[42959]=5998;
squeal_samples[42960]=3414;
squeal_samples[42961]=5215;
squeal_samples[42962]=8035;
squeal_samples[42963]=10747;
squeal_samples[42964]=13335;
squeal_samples[42965]=15806;
squeal_samples[42966]=18171;
squeal_samples[42967]=20425;
squeal_samples[42968]=22589;
squeal_samples[42969]=24648;
squeal_samples[42970]=26627;
squeal_samples[42971]=28508;
squeal_samples[42972]=30305;
squeal_samples[42973]=32025;
squeal_samples[42974]=33668;
squeal_samples[42975]=35237;
squeal_samples[42976]=36734;
squeal_samples[42977]=38167;
squeal_samples[42978]=39528;
squeal_samples[42979]=40836;
squeal_samples[42980]=42078;
squeal_samples[42981]=43272;
squeal_samples[42982]=44406;
squeal_samples[42983]=45490;
squeal_samples[42984]=46528;
squeal_samples[42985]=47515;
squeal_samples[42986]=48460;
squeal_samples[42987]=49361;
squeal_samples[42988]=50224;
squeal_samples[42989]=51043;
squeal_samples[42990]=51834;
squeal_samples[42991]=52581;
squeal_samples[42992]=53303;
squeal_samples[42993]=53986;
squeal_samples[42994]=54645;
squeal_samples[42995]=53929;
squeal_samples[42996]=48334;
squeal_samples[42997]=42628;
squeal_samples[42998]=37289;
squeal_samples[42999]=32295;
squeal_samples[43000]=27618;
squeal_samples[43001]=23237;
squeal_samples[43002]=19139;
squeal_samples[43003]=15306;
squeal_samples[43004]=11724;
squeal_samples[43005]=8358;
squeal_samples[43006]=5226;
squeal_samples[43007]=3410;
squeal_samples[43008]=5920;
squeal_samples[43009]=8719;
squeal_samples[43010]=11393;
squeal_samples[43011]=13954;
squeal_samples[43012]=16403;
squeal_samples[43013]=18731;
squeal_samples[43014]=20968;
squeal_samples[43015]=23103;
squeal_samples[43016]=25145;
squeal_samples[43017]=27094;
squeal_samples[43018]=28954;
squeal_samples[43019]=30734;
squeal_samples[43020]=32434;
squeal_samples[43021]=34053;
squeal_samples[43022]=35609;
squeal_samples[43023]=37086;
squeal_samples[43024]=38505;
squeal_samples[43025]=39849;
squeal_samples[43026]=41140;
squeal_samples[43027]=42374;
squeal_samples[43028]=43547;
squeal_samples[43029]=44674;
squeal_samples[43030]=45742;
squeal_samples[43031]=46766;
squeal_samples[43032]=47746;
squeal_samples[43033]=48675;
squeal_samples[43034]=49575;
squeal_samples[43035]=50420;
squeal_samples[43036]=51236;
squeal_samples[43037]=52013;
squeal_samples[43038]=52756;
squeal_samples[43039]=53466;
squeal_samples[43040]=54140;
squeal_samples[43041]=54793;
squeal_samples[43042]=53485;
squeal_samples[43043]=47661;
squeal_samples[43044]=41998;
squeal_samples[43045]=36699;
squeal_samples[43046]=31741;
squeal_samples[43047]=27098;
squeal_samples[43048]=22751;
squeal_samples[43049]=18680;
squeal_samples[43050]=14883;
squeal_samples[43051]=11318;
squeal_samples[43052]=7989;
squeal_samples[43053]=4871;
squeal_samples[43054]=3574;
squeal_samples[43055]=6303;
squeal_samples[43056]=9077;
squeal_samples[43057]=11742;
squeal_samples[43058]=14283;
squeal_samples[43059]=16714;
squeal_samples[43060]=19036;
squeal_samples[43061]=21252;
squeal_samples[43062]=23378;
squeal_samples[43063]=25406;
squeal_samples[43064]=27343;
squeal_samples[43065]=29196;
squeal_samples[43066]=30962;
squeal_samples[43067]=32652;
squeal_samples[43068]=34260;
squeal_samples[43069]=35806;
squeal_samples[43070]=37270;
squeal_samples[43071]=38682;
squeal_samples[43072]=40022;
squeal_samples[43073]=41305;
squeal_samples[43074]=42525;
squeal_samples[43075]=43697;
squeal_samples[43076]=44808;
squeal_samples[43077]=45880;
squeal_samples[43078]=46892;
squeal_samples[43079]=47865;
squeal_samples[43080]=48792;
squeal_samples[43081]=49679;
squeal_samples[43082]=50522;
squeal_samples[43083]=51337;
squeal_samples[43084]=52104;
squeal_samples[43085]=52846;
squeal_samples[43086]=53549;
squeal_samples[43087]=54222;
squeal_samples[43088]=54872;
squeal_samples[43089]=52870;
squeal_samples[43090]=46929;
squeal_samples[43091]=41316;
squeal_samples[43092]=36058;
squeal_samples[43093]=31141;
squeal_samples[43094]=26533;
squeal_samples[43095]=22224;
squeal_samples[43096]=18189;
squeal_samples[43097]=14421;
squeal_samples[43098]=10885;
squeal_samples[43099]=7579;
squeal_samples[43100]=4482;
squeal_samples[43101]=3808;
squeal_samples[43102]=6648;
squeal_samples[43103]=9412;
squeal_samples[43104]=12058;
squeal_samples[43105]=14586;
squeal_samples[43106]=17006;
squeal_samples[43107]=19311;
squeal_samples[43108]=21516;
squeal_samples[43109]=23628;
squeal_samples[43110]=25645;
squeal_samples[43111]=27573;
squeal_samples[43112]=29413;
squeal_samples[43113]=31169;
squeal_samples[43114]=32850;
squeal_samples[43115]=34449;
squeal_samples[43116]=35988;
squeal_samples[43117]=37444;
squeal_samples[43118]=38845;
squeal_samples[43119]=40175;
squeal_samples[43120]=41453;
squeal_samples[43121]=42667;
squeal_samples[43122]=43829;
squeal_samples[43123]=44939;
squeal_samples[43124]=46000;
squeal_samples[43125]=47006;
squeal_samples[43126]=47977;
squeal_samples[43127]=48894;
squeal_samples[43128]=49784;
squeal_samples[43129]=50616;
squeal_samples[43130]=51424;
squeal_samples[43131]=52193;
squeal_samples[43132]=52929;
squeal_samples[43133]=53623;
squeal_samples[43134]=54299;
squeal_samples[43135]=54939;
squeal_samples[43136]=52149;
squeal_samples[43137]=46192;
squeal_samples[43138]=40629;
squeal_samples[43139]=35413;
squeal_samples[43140]=30537;
squeal_samples[43141]=25973;
squeal_samples[43142]=21691;
squeal_samples[43143]=17692;
squeal_samples[43144]=13954;
squeal_samples[43145]=10452;
squeal_samples[43146]=7171;
squeal_samples[43147]=4105;
squeal_samples[43148]=4117;
squeal_samples[43149]=6988;
squeal_samples[43150]=9738;
squeal_samples[43151]=12374;
squeal_samples[43152]=14887;
squeal_samples[43153]=17283;
squeal_samples[43154]=19584;
squeal_samples[43155]=21777;
squeal_samples[43156]=23879;
squeal_samples[43157]=25879;
squeal_samples[43158]=27798;
squeal_samples[43159]=29624;
squeal_samples[43160]=31373;
squeal_samples[43161]=33043;
squeal_samples[43162]=34639;
squeal_samples[43163]=36157;
squeal_samples[43164]=37613;
squeal_samples[43165]=38999;
squeal_samples[43166]=40331;
squeal_samples[43167]=41594;
squeal_samples[43168]=42804;
squeal_samples[43169]=43959;
squeal_samples[43170]=45061;
squeal_samples[43171]=46119;
squeal_samples[43172]=47123;
squeal_samples[43173]=48084;
squeal_samples[43174]=49000;
squeal_samples[43175]=49877;
squeal_samples[43176]=50709;
squeal_samples[43177]=51513;
squeal_samples[43178]=52274;
squeal_samples[43179]=53007;
squeal_samples[43180]=53703;
squeal_samples[43181]=54366;
squeal_samples[43182]=54957;
squeal_samples[43183]=51367;
squeal_samples[43184]=45470;
squeal_samples[43185]=39949;
squeal_samples[43186]=34779;
squeal_samples[43187]=29941;
squeal_samples[43188]=25408;
squeal_samples[43189]=21172;
squeal_samples[43190]=17203;
squeal_samples[43191]=13495;
squeal_samples[43192]=10018;
squeal_samples[43193]=6769;
squeal_samples[43194]=3771;
squeal_samples[43195]=4468;
squeal_samples[43196]=7336;
squeal_samples[43197]=10062;
squeal_samples[43198]=12687;
squeal_samples[43199]=15179;
squeal_samples[43200]=17568;
squeal_samples[43201]=19849;
squeal_samples[43202]=22036;
squeal_samples[43203]=24122;
squeal_samples[43204]=26116;
squeal_samples[43205]=28019;
squeal_samples[43206]=29838;
squeal_samples[43207]=31574;
squeal_samples[43208]=33234;
squeal_samples[43209]=34820;
squeal_samples[43210]=36336;
squeal_samples[43211]=37783;
squeal_samples[43212]=39162;
squeal_samples[43213]=40485;
squeal_samples[43214]=41740;
squeal_samples[43215]=42942;
squeal_samples[43216]=44089;
squeal_samples[43217]=45187;
squeal_samples[43218]=46235;
squeal_samples[43219]=47237;
squeal_samples[43220]=48190;
squeal_samples[43221]=49103;
squeal_samples[43222]=49974;
squeal_samples[43223]=50806;
squeal_samples[43224]=51597;
squeal_samples[43225]=52362;
squeal_samples[43226]=53079;
squeal_samples[43227]=53783;
squeal_samples[43228]=54438;
squeal_samples[43229]=54860;
squeal_samples[43230]=50597;
squeal_samples[43231]=44754;
squeal_samples[43232]=39270;
squeal_samples[43233]=34147;
squeal_samples[43234]=29342;
squeal_samples[43235]=24858;
squeal_samples[43236]=20648;
squeal_samples[43237]=16726;
squeal_samples[43238]=13035;
squeal_samples[43239]=9592;
squeal_samples[43240]=6369;
squeal_samples[43241]=3529;
squeal_samples[43242]=4829;
squeal_samples[43243]=7667;
squeal_samples[43244]=10395;
squeal_samples[43245]=12987;
squeal_samples[43246]=15478;
squeal_samples[43247]=17848;
squeal_samples[43248]=20119;
squeal_samples[43249]=22290;
squeal_samples[43250]=24368;
squeal_samples[43251]=26350;
squeal_samples[43252]=28243;
squeal_samples[43253]=30051;
squeal_samples[43254]=31775;
squeal_samples[43255]=33432;
squeal_samples[43256]=35003;
squeal_samples[43257]=36513;
squeal_samples[43258]=37951;
squeal_samples[43259]=39321;
squeal_samples[43260]=40633;
squeal_samples[43261]=41881;
squeal_samples[43262]=43079;
squeal_samples[43263]=44221;
squeal_samples[43264]=45314;
squeal_samples[43265]=46352;
squeal_samples[43266]=47350;
squeal_samples[43267]=48295;
squeal_samples[43268]=49206;
squeal_samples[43269]=50067;
squeal_samples[43270]=50897;
squeal_samples[43271]=51689;
squeal_samples[43272]=52437;
squeal_samples[43273]=53170;
squeal_samples[43274]=53850;
squeal_samples[43275]=54512;
squeal_samples[43276]=54662;
squeal_samples[43277]=49834;
squeal_samples[43278]=44040;
squeal_samples[43279]=38602;
squeal_samples[43280]=33524;
squeal_samples[43281]=28758;
squeal_samples[43282]=24303;
squeal_samples[43283]=20131;
squeal_samples[43284]=16233;
squeal_samples[43285]=12586;
squeal_samples[43286]=9165;
squeal_samples[43287]=5971;
squeal_samples[43288]=3382;
squeal_samples[43289]=5182;
squeal_samples[43290]=8009;
squeal_samples[43291]=10712;
squeal_samples[43292]=13301;
squeal_samples[43293]=15770;
squeal_samples[43294]=18127;
squeal_samples[43295]=20386;
squeal_samples[43296]=22545;
squeal_samples[43297]=24610;
squeal_samples[43298]=26575;
squeal_samples[43299]=28466;
squeal_samples[43300]=30258;
squeal_samples[43301]=31982;
squeal_samples[43302]=33620;
squeal_samples[43303]=35184;
squeal_samples[43304]=36683;
squeal_samples[43305]=38112;
squeal_samples[43306]=39477;
squeal_samples[43307]=40784;
squeal_samples[43308]=42024;
squeal_samples[43309]=43215;
squeal_samples[43310]=44352;
squeal_samples[43311]=45434;
squeal_samples[43312]=46470;
squeal_samples[43313]=47456;
squeal_samples[43314]=48401;
squeal_samples[43315]=49305;
squeal_samples[43316]=50163;
squeal_samples[43317]=50990;
squeal_samples[43318]=51770;
squeal_samples[43319]=52528;
squeal_samples[43320]=53240;
squeal_samples[43321]=53926;
squeal_samples[43322]=54583;
squeal_samples[43323]=54352;
squeal_samples[43324]=49083;
squeal_samples[43325]=43327;
squeal_samples[43326]=37936;
squeal_samples[43327]=32900;
squeal_samples[43328]=28174;
squeal_samples[43329]=23759;
squeal_samples[43330]=19624;
squeal_samples[43331]=15754;
squeal_samples[43332]=12137;
squeal_samples[43333]=8743;
squeal_samples[43334]=5574;
squeal_samples[43335]=3330;
squeal_samples[43336]=5529;
squeal_samples[43337]=8343;
squeal_samples[43338]=11027;
squeal_samples[43339]=13608;
squeal_samples[43340]=16057;
squeal_samples[43341]=18406;
squeal_samples[43342]=20652;
squeal_samples[43343]=22803;
squeal_samples[43344]=24846;
squeal_samples[43345]=26810;
squeal_samples[43346]=28677;
squeal_samples[43347]=30473;
squeal_samples[43348]=32177;
squeal_samples[43349]=33810;
squeal_samples[43350]=35366;
squeal_samples[43351]=36860;
squeal_samples[43352]=38275;
squeal_samples[43353]=39635;
squeal_samples[43354]=40932;
squeal_samples[43355]=42165;
squeal_samples[43356]=43353;
squeal_samples[43357]=44477;
squeal_samples[43358]=45560;
squeal_samples[43359]=46582;
squeal_samples[43360]=47570;
squeal_samples[43361]=48502;
squeal_samples[43362]=49410;
squeal_samples[43363]=50256;
squeal_samples[43364]=51082;
squeal_samples[43365]=51854;
squeal_samples[43366]=52610;
squeal_samples[43367]=53317;
squeal_samples[43368]=54001;
squeal_samples[43369]=54652;
squeal_samples[43370]=54415;
squeal_samples[43371]=49146;
squeal_samples[43372]=43386;
squeal_samples[43373]=37992;
squeal_samples[43374]=32945;
squeal_samples[43375]=28215;
squeal_samples[43376]=23802;
squeal_samples[43377]=19659;
squeal_samples[43378]=15791;
squeal_samples[43379]=12168;
squeal_samples[43380]=8772;
squeal_samples[43381]=5601;
squeal_samples[43382]=3354;
squeal_samples[43383]=5552;
squeal_samples[43384]=8363;
squeal_samples[43385]=11053;
squeal_samples[43386]=13622;
squeal_samples[43387]=16077;
squeal_samples[43388]=18421;
squeal_samples[43389]=20670;
squeal_samples[43390]=22814;
squeal_samples[43391]=24865;
squeal_samples[43392]=26825;
squeal_samples[43393]=28691;
squeal_samples[43394]=30482;
squeal_samples[43395]=32186;
squeal_samples[43396]=33819;
squeal_samples[43397]=35375;
squeal_samples[43398]=36865;
squeal_samples[43399]=38281;
squeal_samples[43400]=39644;
squeal_samples[43401]=40934;
squeal_samples[43402]=42175;
squeal_samples[43403]=43352;
squeal_samples[43404]=44479;
squeal_samples[43405]=45561;
squeal_samples[43406]=46583;
squeal_samples[43407]=47570;
squeal_samples[43408]=48504;
squeal_samples[43409]=49405;
squeal_samples[43410]=50258;
squeal_samples[43411]=51076;
squeal_samples[43412]=51857;
squeal_samples[43413]=52603;
squeal_samples[43414]=53314;
squeal_samples[43415]=53998;
squeal_samples[43416]=54650;
squeal_samples[43417]=54414;
squeal_samples[43418]=49138;
squeal_samples[43419]=43384;
squeal_samples[43420]=37987;
squeal_samples[43421]=32939;
squeal_samples[43422]=28214;
squeal_samples[43423]=23794;
squeal_samples[43424]=19652;
squeal_samples[43425]=15785;
squeal_samples[43426]=12157;
squeal_samples[43427]=8771;
squeal_samples[43428]=5593;
squeal_samples[43429]=3352;
squeal_samples[43430]=5546;
squeal_samples[43431]=8360;
squeal_samples[43432]=11042;
squeal_samples[43433]=13614;
squeal_samples[43434]=16070;
squeal_samples[43435]=18418;
squeal_samples[43436]=20661;
squeal_samples[43437]=22802;
squeal_samples[43438]=24858;
squeal_samples[43439]=26813;
squeal_samples[43440]=28687;
squeal_samples[43441]=30473;
squeal_samples[43442]=32180;
squeal_samples[43443]=33810;
squeal_samples[43444]=35366;
squeal_samples[43445]=36854;
squeal_samples[43446]=38272;
squeal_samples[43447]=39632;
squeal_samples[43448]=40926;
squeal_samples[43449]=42165;
squeal_samples[43450]=43348;
squeal_samples[43451]=44473;
squeal_samples[43452]=45552;
squeal_samples[43453]=46579;
squeal_samples[43454]=47564;
squeal_samples[43455]=48502;
squeal_samples[43456]=49398;
squeal_samples[43457]=50250;
squeal_samples[43458]=51071;
squeal_samples[43459]=51847;
squeal_samples[43460]=52593;
squeal_samples[43461]=53304;
squeal_samples[43462]=53989;
squeal_samples[43463]=54639;
squeal_samples[43464]=54405;
squeal_samples[43465]=49128;
squeal_samples[43466]=43374;
squeal_samples[43467]=37977;
squeal_samples[43468]=32935;
squeal_samples[43469]=28203;
squeal_samples[43470]=23786;
squeal_samples[43471]=19640;
squeal_samples[43472]=15777;
squeal_samples[43473]=12147;
squeal_samples[43474]=8759;
squeal_samples[43475]=5586;
squeal_samples[43476]=3339;
squeal_samples[43477]=5539;
squeal_samples[43478]=8349;
squeal_samples[43479]=11032;
squeal_samples[43480]=13603;
squeal_samples[43481]=16063;
squeal_samples[43482]=18406;
squeal_samples[43483]=20653;
squeal_samples[43484]=22791;
squeal_samples[43485]=24848;
squeal_samples[43486]=26803;
squeal_samples[43487]=28679;
squeal_samples[43488]=30460;
squeal_samples[43489]=32175;
squeal_samples[43490]=33796;
squeal_samples[43491]=35359;
squeal_samples[43492]=36840;
squeal_samples[43493]=38267;
squeal_samples[43494]=39619;
squeal_samples[43495]=40919;
squeal_samples[43496]=42152;
squeal_samples[43497]=43340;
squeal_samples[43498]=44462;
squeal_samples[43499]=45544;
squeal_samples[43500]=46567;
squeal_samples[43501]=47556;
squeal_samples[43502]=48490;
squeal_samples[43503]=49391;
squeal_samples[43504]=50237;
squeal_samples[43505]=51064;
squeal_samples[43506]=51834;
squeal_samples[43507]=52586;
squeal_samples[43508]=53293;
squeal_samples[43509]=53980;
squeal_samples[43510]=54627;
squeal_samples[43511]=54397;
squeal_samples[43512]=49116;
squeal_samples[43513]=43367;
squeal_samples[43514]=37965;
squeal_samples[43515]=32926;
squeal_samples[43516]=28193;
squeal_samples[43517]=23775;
squeal_samples[43518]=19633;
squeal_samples[43519]=15763;
squeal_samples[43520]=12141;
squeal_samples[43521]=8747;
squeal_samples[43522]=5577;
squeal_samples[43523]=3330;
squeal_samples[43524]=5528;
squeal_samples[43525]=8339;
squeal_samples[43526]=11023;
squeal_samples[43527]=13593;
squeal_samples[43528]=16052;
squeal_samples[43529]=18399;
squeal_samples[43530]=20639;
squeal_samples[43531]=22785;
squeal_samples[43532]=24835;
squeal_samples[43533]=26796;
squeal_samples[43534]=28666;
squeal_samples[43535]=30454;
squeal_samples[43536]=32160;
squeal_samples[43537]=33791;
squeal_samples[43538]=35345;
squeal_samples[43539]=36835;
squeal_samples[43540]=38253;
squeal_samples[43541]=39611;
squeal_samples[43542]=40908;
squeal_samples[43543]=42144;
squeal_samples[43544]=43328;
squeal_samples[43545]=44456;
squeal_samples[43546]=45528;
squeal_samples[43547]=46564;
squeal_samples[43548]=47541;
squeal_samples[43549]=48483;
squeal_samples[43550]=49379;
squeal_samples[43551]=50229;
squeal_samples[43552]=51053;
squeal_samples[43553]=51826;
squeal_samples[43554]=52573;
squeal_samples[43555]=53286;
squeal_samples[43556]=53966;
squeal_samples[43557]=54623;
squeal_samples[43558]=54382;
squeal_samples[43559]=49111;
squeal_samples[43560]=43352;
squeal_samples[43561]=37959;
squeal_samples[43562]=32914;
squeal_samples[43563]=28184;
squeal_samples[43564]=23766;
squeal_samples[43565]=19620;
squeal_samples[43566]=15759;
squeal_samples[43567]=12125;
squeal_samples[43568]=8742;
squeal_samples[43569]=5563;
squeal_samples[43570]=3323;
squeal_samples[43571]=5517;
squeal_samples[43572]=8330;
squeal_samples[43573]=11013;
squeal_samples[43574]=13581;
squeal_samples[43575]=16046;
squeal_samples[43576]=18385;
squeal_samples[43577]=20633;
squeal_samples[43578]=22772;
squeal_samples[43579]=24827;
squeal_samples[43580]=26785;
squeal_samples[43581]=28658;
squeal_samples[43582]=30442;
squeal_samples[43583]=32152;
squeal_samples[43584]=33779;
squeal_samples[43585]=35338;
squeal_samples[43586]=36822;
squeal_samples[43587]=38246;
squeal_samples[43588]=39600;
squeal_samples[43589]=40897;
squeal_samples[43590]=42136;
squeal_samples[43591]=43317;
squeal_samples[43592]=44445;
squeal_samples[43593]=45522;
squeal_samples[43594]=46550;
squeal_samples[43595]=47533;
squeal_samples[43596]=48474;
squeal_samples[43597]=49368;
squeal_samples[43598]=50219;
squeal_samples[43599]=51045;
squeal_samples[43600]=51814;
squeal_samples[43601]=52564;
squeal_samples[43602]=53278;
squeal_samples[43603]=53954;
squeal_samples[43604]=54615;
squeal_samples[43605]=54372;
squeal_samples[43606]=49099;
squeal_samples[43607]=43345;
squeal_samples[43608]=37948;
squeal_samples[43609]=32905;
squeal_samples[43610]=28173;
squeal_samples[43611]=23758;
squeal_samples[43612]=19608;
squeal_samples[43613]=15751;
squeal_samples[43614]=12114;
squeal_samples[43615]=8732;
squeal_samples[43616]=5555;
squeal_samples[43617]=3311;
squeal_samples[43618]=5509;
squeal_samples[43619]=8319;
squeal_samples[43620]=11003;
squeal_samples[43621]=13574;
squeal_samples[43622]=16031;
squeal_samples[43623]=18381;
squeal_samples[43624]=20618;
squeal_samples[43625]=22766;
squeal_samples[43626]=24815;
squeal_samples[43627]=26777;
squeal_samples[43628]=28646;
squeal_samples[43629]=30435;
squeal_samples[43630]=32139;
squeal_samples[43631]=33771;
squeal_samples[43632]=35327;
squeal_samples[43633]=36813;
squeal_samples[43634]=38236;
squeal_samples[43635]=39590;
squeal_samples[43636]=40888;
squeal_samples[43637]=42124;
squeal_samples[43638]=43308;
squeal_samples[43639]=44437;
squeal_samples[43640]=45509;
squeal_samples[43641]=46543;
squeal_samples[43642]=47521;
squeal_samples[43643]=48466;
squeal_samples[43644]=49355;
squeal_samples[43645]=50214;
squeal_samples[43646]=51029;
squeal_samples[43647]=51809;
squeal_samples[43648]=52553;
squeal_samples[43649]=53266;
squeal_samples[43650]=53947;
squeal_samples[43651]=54602;
squeal_samples[43652]=54364;
squeal_samples[43653]=49089;
squeal_samples[43654]=43335;
squeal_samples[43655]=37937;
squeal_samples[43656]=32897;
squeal_samples[43657]=28162;
squeal_samples[43658]=23748;
squeal_samples[43659]=19598;
squeal_samples[43660]=15741;
squeal_samples[43661]=12105;
squeal_samples[43662]=8723;
squeal_samples[43663]=5543;
squeal_samples[43664]=3303;
squeal_samples[43665]=5497;
squeal_samples[43666]=8311;
squeal_samples[43667]=10994;
squeal_samples[43668]=13561;
squeal_samples[43669]=16025;
squeal_samples[43670]=18367;
squeal_samples[43671]=20612;
squeal_samples[43672]=22754;
squeal_samples[43673]=24806;
squeal_samples[43674]=26766;
squeal_samples[43675]=28637;
squeal_samples[43676]=30425;
squeal_samples[43677]=32129;
squeal_samples[43678]=33763;
squeal_samples[43679]=35314;
squeal_samples[43680]=36806;
squeal_samples[43681]=38223;
squeal_samples[43682]=39583;
squeal_samples[43683]=40876;
squeal_samples[43684]=42117;
squeal_samples[43685]=43295;
squeal_samples[43686]=44428;
squeal_samples[43687]=45499;
squeal_samples[43688]=46532;
squeal_samples[43689]=47515;
squeal_samples[43690]=48450;
squeal_samples[43691]=49351;
squeal_samples[43692]=50199;
squeal_samples[43693]=51022;
squeal_samples[43694]=51798;
squeal_samples[43695]=52542;
squeal_samples[43696]=53258;
squeal_samples[43697]=53934;
squeal_samples[43698]=54594;
squeal_samples[43699]=54726;
squeal_samples[43700]=49903;
squeal_samples[43701]=44087;
squeal_samples[43702]=38647;
squeal_samples[43703]=33552;
squeal_samples[43704]=28785;
squeal_samples[43705]=24322;
squeal_samples[43706]=20145;
squeal_samples[43707]=16242;
squeal_samples[43708]=12583;
squeal_samples[43709]=9161;
squeal_samples[43710]=5953;
squeal_samples[43711]=3368;
squeal_samples[43712]=5162;
squeal_samples[43713]=7984;
squeal_samples[43714]=10686;
squeal_samples[43715]=13269;
squeal_samples[43716]=15743;
squeal_samples[43717]=18091;
squeal_samples[43718]=20353;
squeal_samples[43719]=22504;
squeal_samples[43720]=24569;
squeal_samples[43721]=26538;
squeal_samples[43722]=28417;
squeal_samples[43723]=30211;
squeal_samples[43724]=31934;
squeal_samples[43725]=33569;
squeal_samples[43726]=35134;
squeal_samples[43727]=36632;
squeal_samples[43728]=38056;
squeal_samples[43729]=39421;
squeal_samples[43730]=40720;
squeal_samples[43731]=41971;
squeal_samples[43732]=43151;
squeal_samples[43733]=44286;
squeal_samples[43734]=45373;
squeal_samples[43735]=46404;
squeal_samples[43736]=47399;
squeal_samples[43737]=48332;
squeal_samples[43738]=49236;
squeal_samples[43739]=50100;
squeal_samples[43740]=50916;
squeal_samples[43741]=51704;
squeal_samples[43742]=52449;
squeal_samples[43743]=53172;
squeal_samples[43744]=53849;
squeal_samples[43745]=54506;
squeal_samples[43746]=54917;
squeal_samples[43747]=50649;
squeal_samples[43748]=44788;
squeal_samples[43749]=39308;
squeal_samples[43750]=34162;
squeal_samples[43751]=29366;
squeal_samples[43752]=24856;
squeal_samples[43753]=20650;
squeal_samples[43754]=16708;
squeal_samples[43755]=13024;
squeal_samples[43756]=9568;
squeal_samples[43757]=6342;
squeal_samples[43758]=3499;
squeal_samples[43759]=4792;
squeal_samples[43760]=7634;
squeal_samples[43761]=10346;
squeal_samples[43762]=12949;
squeal_samples[43763]=15426;
squeal_samples[43764]=17800;
squeal_samples[43765]=20071;
squeal_samples[43766]=22233;
squeal_samples[43767]=24312;
squeal_samples[43768]=26288;
squeal_samples[43769]=28179;
squeal_samples[43770]=29985;
squeal_samples[43771]=31711;
squeal_samples[43772]=33361;
squeal_samples[43773]=34932;
squeal_samples[43774]=36439;
squeal_samples[43775]=37872;
squeal_samples[43776]=39249;
squeal_samples[43777]=40553;
squeal_samples[43778]=41808;
squeal_samples[43779]=43002;
squeal_samples[43780]=44139;
squeal_samples[43781]=45233;
squeal_samples[43782]=46266;
squeal_samples[43783]=47262;
squeal_samples[43784]=48210;
squeal_samples[43785]=49116;
squeal_samples[43786]=49983;
squeal_samples[43787]=50802;
squeal_samples[43788]=51603;
squeal_samples[43789]=52346;
squeal_samples[43790]=53074;
squeal_samples[43791]=53759;
squeal_samples[43792]=54418;
squeal_samples[43793]=54997;
squeal_samples[43794]=51395;
squeal_samples[43795]=45496;
squeal_samples[43796]=39952;
squeal_samples[43797]=34787;
squeal_samples[43798]=29928;
squeal_samples[43799]=25402;
squeal_samples[43800]=21145;
squeal_samples[43801]=17174;
squeal_samples[43802]=13458;
squeal_samples[43803]=9977;
squeal_samples[43804]=6723;
squeal_samples[43805]=3717;
squeal_samples[43806]=4419;
squeal_samples[43807]=7275;
squeal_samples[43808]=10001;
squeal_samples[43809]=12618;
squeal_samples[43810]=15110;
squeal_samples[43811]=17501;
squeal_samples[43812]=19775;
squeal_samples[43813]=21961;
squeal_samples[43814]=24045;
squeal_samples[43815]=26034;
squeal_samples[43816]=27936;
squeal_samples[43817]=29754;
squeal_samples[43818]=31488;
squeal_samples[43819]=33151;
squeal_samples[43820]=34733;
squeal_samples[43821]=36243;
squeal_samples[43822]=37691;
squeal_samples[43823]=39069;
squeal_samples[43824]=40387;
squeal_samples[43825]=41640;
squeal_samples[43826]=42847;
squeal_samples[43827]=43986;
squeal_samples[43828]=45090;
squeal_samples[43829]=46129;
squeal_samples[43830]=47135;
squeal_samples[43831]=48085;
squeal_samples[43832]=48998;
squeal_samples[43833]=49869;
squeal_samples[43834]=50696;
squeal_samples[43835]=51493;
squeal_samples[43836]=52246;
squeal_samples[43837]=52977;
squeal_samples[43838]=53665;
squeal_samples[43839]=54331;
squeal_samples[43840]=54958;
squeal_samples[43841]=52164;
squeal_samples[43842]=46196;
squeal_samples[43843]=40624;
squeal_samples[43844]=35400;
squeal_samples[43845]=30515;
squeal_samples[43846]=25937;
squeal_samples[43847]=21653;
squeal_samples[43848]=17647;
squeal_samples[43849]=13900;
squeal_samples[43850]=10389;
squeal_samples[43851]=7112;
squeal_samples[43852]=4031;
squeal_samples[43853]=4041;
squeal_samples[43854]=6912;
squeal_samples[43855]=9659;
squeal_samples[43856]=12288;
squeal_samples[43857]=14797;
squeal_samples[43858]=17196;
squeal_samples[43859]=19490;
squeal_samples[43860]=21684;
squeal_samples[43861]=23781;
squeal_samples[43862]=25780;
squeal_samples[43863]=27698;
squeal_samples[43864]=29521;
squeal_samples[43865]=31267;
squeal_samples[43866]=32936;
squeal_samples[43867]=34527;
squeal_samples[43868]=36049;
squeal_samples[43869]=37501;
squeal_samples[43870]=38893;
squeal_samples[43871]=40212;
squeal_samples[43872]=41481;
squeal_samples[43873]=42687;
squeal_samples[43874]=43840;
squeal_samples[43875]=44939;
squeal_samples[43876]=45995;
squeal_samples[43877]=46994;
squeal_samples[43878]=47961;
squeal_samples[43879]=48871;
squeal_samples[43880]=49752;
squeal_samples[43881]=50582;
squeal_samples[43882]=51388;
squeal_samples[43883]=52141;
squeal_samples[43884]=52876;
squeal_samples[43885]=53569;
squeal_samples[43886]=54235;
squeal_samples[43887]=54878;
squeal_samples[43888]=52866;
squeal_samples[43889]=46913;
squeal_samples[43890]=41290;
squeal_samples[43891]=36026;
squeal_samples[43892]=31098;
squeal_samples[43893]=26481;
squeal_samples[43894]=22164;
squeal_samples[43895]=18127;
squeal_samples[43896]=14343;
squeal_samples[43897]=10813;
squeal_samples[43898]=7494;
squeal_samples[43899]=4402;
squeal_samples[43900]=3706;
squeal_samples[43901]=6556;
squeal_samples[43902]=9313;
squeal_samples[43903]=11954;
squeal_samples[43904]=14483;
squeal_samples[43905]=16893;
squeal_samples[43906]=19203;
squeal_samples[43907]=21400;
squeal_samples[43908]=23516;
squeal_samples[43909]=25527;
squeal_samples[43910]=27448;
squeal_samples[43911]=29289;
squeal_samples[43912]=31048;
squeal_samples[43913]=32721;
squeal_samples[43914]=34327;
squeal_samples[43915]=35851;
squeal_samples[43916]=37314;
squeal_samples[43917]=38709;
squeal_samples[43918]=40040;
squeal_samples[43919]=41319;
squeal_samples[43920]=42526;
squeal_samples[43921]=43688;
squeal_samples[43922]=44800;
squeal_samples[43923]=45860;
squeal_samples[43924]=46865;
squeal_samples[43925]=47836;
squeal_samples[43926]=48750;
squeal_samples[43927]=49630;
squeal_samples[43928]=50474;
squeal_samples[43929]=51275;
squeal_samples[43930]=52042;
squeal_samples[43931]=52778;
squeal_samples[43932]=53473;
squeal_samples[43933]=54143;
squeal_samples[43934]=54786;
squeal_samples[43935]=53470;
squeal_samples[43936]=47632;
squeal_samples[43937]=41964;
squeal_samples[43938]=36652;
squeal_samples[43939]=31686;
squeal_samples[43940]=27028;
squeal_samples[43941]=22685;
squeal_samples[43942]=18602;
squeal_samples[43943]=14797;
squeal_samples[43944]=11232;
squeal_samples[43945]=7886;
squeal_samples[43946]=4767;
squeal_samples[43947]=3469;
squeal_samples[43948]=6189;
squeal_samples[43949]=8970;
squeal_samples[43950]=11624;
squeal_samples[43951]=14160;
squeal_samples[43952]=16591;
squeal_samples[43953]=18903;
squeal_samples[43954]=21130;
squeal_samples[43955]=23244;
squeal_samples[43956]=25266;
squeal_samples[43957]=27209;
squeal_samples[43958]=29054;
squeal_samples[43959]=30820;
squeal_samples[43960]=32509;
squeal_samples[43961]=34117;
squeal_samples[43962]=35655;
squeal_samples[43963]=37125;
squeal_samples[43964]=38529;
squeal_samples[43965]=39869;
squeal_samples[43966]=41152;
squeal_samples[43967]=42369;
squeal_samples[43968]=43538;
squeal_samples[43969]=44655;
squeal_samples[43970]=45718;
squeal_samples[43971]=46733;
squeal_samples[43972]=47706;
squeal_samples[43973]=48630;
squeal_samples[43974]=49521;
squeal_samples[43975]=50356;
squeal_samples[43976]=51172;
squeal_samples[43977]=51937;
squeal_samples[43978]=52677;
squeal_samples[43979]=53380;
squeal_samples[43980]=54054;
squeal_samples[43981]=54697;
squeal_samples[43982]=53973;
squeal_samples[43983]=48360;
squeal_samples[43984]=42638;
squeal_samples[43985]=37291;
squeal_samples[43986]=32275;
squeal_samples[43987]=27594;
squeal_samples[43988]=23195;
squeal_samples[43989]=19092;
squeal_samples[43990]=15247;
squeal_samples[43991]=11649;
squeal_samples[43992]=8282;
squeal_samples[43993]=5134;
squeal_samples[43994]=3320;
squeal_samples[43995]=5822;
squeal_samples[43996]=8614;
squeal_samples[43997]=11291;
squeal_samples[43998]=13840;
squeal_samples[43999]=16287;
squeal_samples[44000]=18613;
squeal_samples[44001]=20848;
squeal_samples[44002]=22972;
squeal_samples[44003]=25016;
squeal_samples[44004]=26956;
squeal_samples[44005]=28818;
squeal_samples[44006]=30596;
squeal_samples[44007]=32287;
squeal_samples[44008]=33914;
squeal_samples[44009]=35454;
squeal_samples[44010]=36940;
squeal_samples[44011]=38344;
squeal_samples[44012]=39699;
squeal_samples[44013]=40981;
squeal_samples[44014]=42211;
squeal_samples[44015]=43384;
squeal_samples[44016]=44507;
squeal_samples[44017]=45576;
squeal_samples[44018]=46600;
squeal_samples[44019]=47575;
squeal_samples[44020]=48509;
squeal_samples[44021]=49399;
squeal_samples[44022]=50247;
squeal_samples[44023]=51061;
squeal_samples[44024]=51833;
squeal_samples[44025]=52578;
squeal_samples[44026]=53283;
squeal_samples[44027]=53963;
squeal_samples[44028]=54610;
squeal_samples[44029]=54367;
squeal_samples[44030]=49087;
squeal_samples[44031]=43326;
squeal_samples[44032]=37930;
squeal_samples[44033]=32876;
squeal_samples[44034]=28147;
squeal_samples[44035]=23719;
squeal_samples[44036]=19580;
squeal_samples[44037]=15706;
squeal_samples[44038]=12078;
squeal_samples[44039]=8686;
squeal_samples[44040]=5504;
squeal_samples[44041]=3262;
squeal_samples[44042]=5452;
squeal_samples[44043]=8264;
squeal_samples[44044]=10947;
squeal_samples[44045]=13518;
squeal_samples[44046]=15976;
squeal_samples[44047]=18319;
squeal_samples[44048]=20558;
squeal_samples[44049]=22704;
squeal_samples[44050]=24754;
squeal_samples[44051]=26710;
squeal_samples[44052]=28579;
squeal_samples[44053]=30370;
squeal_samples[44054]=32065;
squeal_samples[44055]=33709;
squeal_samples[44056]=35254;
squeal_samples[44057]=36753;
squeal_samples[44058]=38158;
squeal_samples[44059]=39521;
squeal_samples[44060]=40817;
squeal_samples[44061]=42050;
squeal_samples[44062]=43234;
squeal_samples[44063]=44354;
squeal_samples[44064]=45442;
squeal_samples[44065]=46462;
squeal_samples[44066]=47446;
squeal_samples[44067]=48387;
squeal_samples[44068]=49278;
squeal_samples[44069]=50136;
squeal_samples[44070]=50947;
squeal_samples[44071]=51729;
squeal_samples[44072]=52477;
squeal_samples[44073]=53187;
squeal_samples[44074]=53869;
squeal_samples[44075]=54519;
squeal_samples[44076]=54924;
squeal_samples[44077]=50656;
squeal_samples[44078]=44786;
squeal_samples[44079]=39297;
squeal_samples[44080]=34156;
squeal_samples[44081]=29349;
squeal_samples[44082]=24839;
squeal_samples[44083]=20628;
squeal_samples[44084]=16684;
squeal_samples[44085]=12993;
squeal_samples[44086]=9538;
squeal_samples[44087]=6307;
squeal_samples[44088]=3460;
squeal_samples[44089]=4759;
squeal_samples[44090]=7595;
squeal_samples[44091]=10309;
squeal_samples[44092]=12904;
squeal_samples[44093]=15386;
squeal_samples[44094]=17753;
squeal_samples[44095]=20024;
squeal_samples[44096]=22194;
squeal_samples[44097]=24262;
squeal_samples[44098]=26243;
squeal_samples[44099]=28132;
squeal_samples[44100]=29939;
squeal_samples[44101]=31663;
squeal_samples[44102]=33309;
squeal_samples[44103]=34881;
squeal_samples[44104]=36385;
squeal_samples[44105]=37822;
squeal_samples[44106]=39195;
squeal_samples[44107]=40501;
squeal_samples[44108]=41751;
squeal_samples[44109]=42943;
squeal_samples[44110]=44083;
squeal_samples[44111]=45174;
squeal_samples[44112]=46214;
squeal_samples[44113]=47205;
squeal_samples[44114]=48150;
squeal_samples[44115]=49063;
squeal_samples[44116]=49918;
squeal_samples[44117]=50753;
squeal_samples[44118]=51530;
squeal_samples[44119]=52298;
squeal_samples[44120]=53003;
squeal_samples[44121]=53707;
squeal_samples[44122]=54350;
squeal_samples[44123]=54989;
squeal_samples[44124]=52175;
squeal_samples[44125]=46219;
squeal_samples[44126]=40631;
squeal_samples[44127]=35409;
squeal_samples[44128]=30515;
squeal_samples[44129]=25933;
squeal_samples[44130]=21649;
squeal_samples[44131]=17637;
squeal_samples[44132]=13888;
squeal_samples[44133]=10377;
squeal_samples[44134]=7089;
squeal_samples[44135]=4013;
squeal_samples[44136]=4018;
squeal_samples[44137]=6891;
squeal_samples[44138]=9635;
squeal_samples[44139]=12260;
squeal_samples[44140]=14766;
squeal_samples[44141]=17167;
squeal_samples[44142]=19454;
squeal_samples[44143]=21658;
squeal_samples[44144]=23743;
squeal_samples[44145]=25748;
squeal_samples[44146]=27660;
squeal_samples[44147]=29484;
squeal_samples[44148]=31231;
squeal_samples[44149]=32896;
squeal_samples[44150]=34489;
squeal_samples[44151]=36008;
squeal_samples[44152]=37463;
squeal_samples[44153]=38846;
squeal_samples[44154]=40175;
squeal_samples[44155]=41435;
squeal_samples[44156]=42641;
squeal_samples[44157]=43797;
squeal_samples[44158]=44896;
squeal_samples[44159]=45954;
squeal_samples[44160]=46951;
squeal_samples[44161]=47913;
squeal_samples[44162]=48824;
squeal_samples[44163]=49703;
squeal_samples[44164]=50536;
squeal_samples[44165]=51337;
squeal_samples[44166]=52096;
squeal_samples[44167]=52826;
squeal_samples[44168]=53522;
squeal_samples[44169]=54188;
squeal_samples[44170]=54821;
squeal_samples[44171]=53506;
squeal_samples[44172]=47656;
squeal_samples[44173]=41988;
squeal_samples[44174]=36667;
squeal_samples[44175]=31703;
squeal_samples[44176]=27039;
squeal_samples[44177]=22690;
squeal_samples[44178]=18601;
squeal_samples[44179]=14799;
squeal_samples[44180]=11225;
squeal_samples[44181]=7881;
squeal_samples[44182]=4757;
squeal_samples[44183]=3456;
squeal_samples[44184]=6176;
squeal_samples[44185]=8952;
squeal_samples[44186]=11601;
squeal_samples[44187]=14148;
squeal_samples[44188]=16568;
squeal_samples[44189]=18889;
squeal_samples[44190]=21103;
squeal_samples[44191]=23224;
squeal_samples[44192]=25246;
squeal_samples[44193]=27179;
squeal_samples[44194]=29029;
squeal_samples[44195]=30793;
squeal_samples[44196]=32481;
squeal_samples[44197]=34085;
squeal_samples[44198]=35628;
squeal_samples[44199]=37092;
squeal_samples[44200]=38497;
squeal_samples[44201]=39837;
squeal_samples[44202]=41119;
squeal_samples[44203]=42336;
squeal_samples[44204]=43506;
squeal_samples[44205]=44617;
squeal_samples[44206]=45679;
squeal_samples[44207]=46698;
squeal_samples[44208]=47663;
squeal_samples[44209]=48598;
squeal_samples[44210]=49477;
squeal_samples[44211]=50323;
squeal_samples[44212]=51130;
squeal_samples[44213]=51902;
squeal_samples[44214]=52637;
squeal_samples[44215]=53338;
squeal_samples[44216]=54013;
squeal_samples[44217]=54660;
squeal_samples[44218]=54412;
squeal_samples[44219]=49128;
squeal_samples[44220]=43354;
squeal_samples[44221]=37958;
squeal_samples[44222]=32901;
squeal_samples[44223]=28168;
squeal_samples[44224]=23735;
squeal_samples[44225]=19595;
squeal_samples[44226]=15714;
squeal_samples[44227]=12086;
squeal_samples[44228]=8687;
squeal_samples[44229]=5506;
squeal_samples[44230]=3258;
squeal_samples[44231]=5452;
squeal_samples[44232]=8258;
squeal_samples[44233]=10940;
squeal_samples[44234]=13513;
squeal_samples[44235]=15963;
squeal_samples[44236]=18306;
squeal_samples[44237]=20548;
squeal_samples[44238]=22690;
squeal_samples[44239]=24740;
squeal_samples[44240]=26696;
squeal_samples[44241]=28563;
squeal_samples[44242]=30350;
squeal_samples[44243]=32053;
squeal_samples[44244]=33679;
squeal_samples[44245]=35240;
squeal_samples[44246]=36722;
squeal_samples[44247]=38142;
squeal_samples[44248]=39495;
squeal_samples[44249]=40794;
squeal_samples[44250]=42024;
squeal_samples[44251]=43208;
squeal_samples[44252]=44336;
squeal_samples[44253]=45410;
squeal_samples[44254]=46436;
squeal_samples[44255]=47418;
squeal_samples[44256]=48357;
squeal_samples[44257]=49253;
squeal_samples[44258]=50104;
squeal_samples[44259]=50922;
squeal_samples[44260]=51700;
squeal_samples[44261]=52451;
squeal_samples[44262]=53149;
squeal_samples[44263]=53841;
squeal_samples[44264]=54485;
squeal_samples[44265]=54902;
squeal_samples[44266]=50619;
squeal_samples[44267]=44754;
squeal_samples[44268]=39267;
squeal_samples[44269]=34125;
squeal_samples[44270]=29314;
squeal_samples[44271]=24807;
squeal_samples[44272]=20593;
squeal_samples[44273]=16652;
squeal_samples[44274]=12959;
squeal_samples[44275]=9506;
squeal_samples[44276]=6270;
squeal_samples[44277]=3431;
squeal_samples[44278]=4717;
squeal_samples[44279]=7559;
squeal_samples[44280]=10273;
squeal_samples[44281]=12871;
squeal_samples[44282]=15354;
squeal_samples[44283]=17719;
squeal_samples[44284]=19990;
squeal_samples[44285]=22155;
squeal_samples[44286]=24228;
squeal_samples[44287]=26206;
squeal_samples[44288]=28092;
squeal_samples[44289]=29900;
squeal_samples[44290]=31626;
squeal_samples[44291]=33273;
squeal_samples[44292]=34850;
squeal_samples[44293]=36350;
squeal_samples[44294]=37783;
squeal_samples[44295]=39158;
squeal_samples[44296]=40461;
squeal_samples[44297]=41719;
squeal_samples[44298]=42908;
squeal_samples[44299]=44051;
squeal_samples[44300]=45134;
squeal_samples[44301]=46177;
squeal_samples[44302]=47170;
squeal_samples[44303]=48113;
squeal_samples[44304]=49021;
squeal_samples[44305]=49885;
squeal_samples[44306]=50707;
squeal_samples[44307]=51500;
squeal_samples[44308]=52249;
squeal_samples[44309]=52973;
squeal_samples[44310]=53661;
squeal_samples[44311]=54319;
squeal_samples[44312]=54943;
squeal_samples[44313]=52142;
squeal_samples[44314]=46175;
squeal_samples[44315]=40596;
squeal_samples[44316]=35369;
squeal_samples[44317]=30477;
squeal_samples[44318]=25898;
squeal_samples[44319]=21612;
squeal_samples[44320]=17597;
squeal_samples[44321]=13850;
squeal_samples[44322]=10340;
squeal_samples[44323]=7046;
squeal_samples[44324]=3978;
squeal_samples[44325]=3976;
squeal_samples[44326]=6857;
squeal_samples[44327]=9592;
squeal_samples[44328]=12223;
squeal_samples[44329]=14733;
squeal_samples[44330]=17124;
squeal_samples[44331]=19423;
squeal_samples[44332]=21612;
squeal_samples[44333]=23709;
squeal_samples[44334]=25712;
squeal_samples[44335]=27621;
squeal_samples[44336]=29446;
squeal_samples[44337]=31192;
squeal_samples[44338]=32858;
squeal_samples[44339]=34448;
squeal_samples[44340]=35972;
squeal_samples[44341]=37421;
squeal_samples[44342]=38812;
squeal_samples[44343]=40130;
squeal_samples[44344]=41401;
squeal_samples[44345]=42599;
squeal_samples[44346]=43760;
squeal_samples[44347]=44859;
squeal_samples[44348]=45912;
squeal_samples[44349]=46914;
squeal_samples[44350]=47873;
squeal_samples[44351]=48787;
squeal_samples[44352]=49663;
squeal_samples[44353]=50500;
squeal_samples[44354]=51294;
squeal_samples[44355]=52062;
squeal_samples[44356]=52783;
squeal_samples[44357]=53487;
squeal_samples[44358]=54147;
squeal_samples[44359]=54782;
squeal_samples[44360]=53469;
squeal_samples[44361]=47616;
squeal_samples[44362]=41950;
squeal_samples[44363]=36629;
squeal_samples[44364]=31662;
squeal_samples[44365]=27002;
squeal_samples[44366]=22650;
squeal_samples[44367]=18569;
squeal_samples[44368]=14761;
squeal_samples[44369]=11183;
squeal_samples[44370]=7848;
squeal_samples[44371]=4711;
squeal_samples[44372]=3424;
squeal_samples[44373]=6133;
squeal_samples[44374]=8914;
squeal_samples[44375]=11564;
squeal_samples[44376]=14107;
squeal_samples[44377]=16531;
squeal_samples[44378]=18850;
squeal_samples[44379]=21062;
squeal_samples[44380]=23189;
squeal_samples[44381]=25204;
squeal_samples[44382]=27142;
squeal_samples[44383]=28989;
squeal_samples[44384]=30756;
squeal_samples[44385]=32439;
squeal_samples[44386]=34050;
squeal_samples[44387]=35587;
squeal_samples[44388]=37053;
squeal_samples[44389]=38460;
squeal_samples[44390]=39796;
squeal_samples[44391]=41081;
squeal_samples[44392]=42298;
squeal_samples[44393]=43466;
squeal_samples[44394]=44579;
squeal_samples[44395]=45641;
squeal_samples[44396]=46657;
squeal_samples[44397]=47627;
squeal_samples[44398]=48556;
squeal_samples[44399]=49441;
squeal_samples[44400]=50283;
squeal_samples[44401]=51090;
squeal_samples[44402]=51866;
squeal_samples[44403]=52594;
squeal_samples[44404]=53302;
squeal_samples[44405]=53973;
squeal_samples[44406]=54620;
squeal_samples[44407]=54749;
squeal_samples[44408]=49908;
squeal_samples[44409]=44088;
squeal_samples[44410]=38636;
squeal_samples[44411]=33535;
squeal_samples[44412]=28759;
squeal_samples[44413]=24288;
squeal_samples[44414]=20105;
squeal_samples[44415]=16192;
squeal_samples[44416]=12528;
squeal_samples[44417]=9102;
squeal_samples[44418]=5888;
squeal_samples[44419]=3298;
squeal_samples[44420]=5086;
squeal_samples[44421]=7909;
squeal_samples[44422]=10603;
squeal_samples[44423]=13186;
squeal_samples[44424]=15652;
squeal_samples[44425]=18009;
squeal_samples[44426]=20257;
squeal_samples[44427]=22414;
squeal_samples[44428]=24473;
squeal_samples[44429]=26434;
squeal_samples[44430]=28319;
squeal_samples[44431]=30111;
squeal_samples[44432]=31822;
squeal_samples[44433]=33464;
squeal_samples[44434]=35025;
squeal_samples[44435]=36517;
squeal_samples[44436]=37944;
squeal_samples[44437]=39307;
squeal_samples[44438]=40606;
squeal_samples[44439]=41853;
squeal_samples[44440]=43035;
squeal_samples[44441]=44170;
squeal_samples[44442]=45250;
squeal_samples[44443]=46284;
squeal_samples[44444]=47271;
squeal_samples[44445]=48214;
squeal_samples[44446]=49112;
squeal_samples[44447]=49968;
squeal_samples[44448]=50789;
squeal_samples[44449]=51576;
squeal_samples[44450]=52321;
squeal_samples[44451]=53041;
squeal_samples[44452]=53716;
squeal_samples[44453]=54379;
squeal_samples[44454]=55000;
squeal_samples[44455]=52194;
squeal_samples[44456]=46218;
squeal_samples[44457]=40636;
squeal_samples[44458]=35404;
squeal_samples[44459]=30509;
squeal_samples[44460]=25923;
squeal_samples[44461]=21636;
squeal_samples[44462]=17619;
squeal_samples[44463]=13868;
squeal_samples[44464]=10354;
squeal_samples[44465]=7062;
squeal_samples[44466]=3986;
squeal_samples[44467]=3986;
squeal_samples[44468]=6858;
squeal_samples[44469]=9598;
squeal_samples[44470]=12225;
squeal_samples[44471]=14733;
squeal_samples[44472]=17127;
squeal_samples[44473]=19419;
squeal_samples[44474]=21612;
squeal_samples[44475]=23702;
squeal_samples[44476]=25704;
squeal_samples[44477]=27614;
squeal_samples[44478]=29438;
squeal_samples[44479]=31185;
squeal_samples[44480]=32851;
squeal_samples[44481]=34441;
squeal_samples[44482]=35958;
squeal_samples[44483]=37409;
squeal_samples[44484]=38797;
squeal_samples[44485]=40121;
squeal_samples[44486]=41385;
squeal_samples[44487]=42588;
squeal_samples[44488]=43746;
squeal_samples[44489]=44841;
squeal_samples[44490]=45892;
squeal_samples[44491]=46900;
squeal_samples[44492]=47855;
squeal_samples[44493]=48774;
squeal_samples[44494]=49640;
squeal_samples[44495]=50483;
squeal_samples[44496]=51277;
squeal_samples[44497]=52041;
squeal_samples[44498]=52763;
squeal_samples[44499]=53459;
squeal_samples[44500]=54124;
squeal_samples[44501]=54766;
squeal_samples[44502]=54027;
squeal_samples[44503]=48406;
squeal_samples[44504]=42679;
squeal_samples[44505]=37311;
squeal_samples[44506]=32297;
squeal_samples[44507]=27597;
squeal_samples[44508]=23200;
squeal_samples[44509]=19086;
squeal_samples[44510]=15238;
squeal_samples[44511]=11636;
squeal_samples[44512]=8261;
squeal_samples[44513]=5103;
squeal_samples[44514]=3291;
squeal_samples[44515]=5781;
squeal_samples[44516]=8578;
squeal_samples[44517]=11239;
squeal_samples[44518]=13797;
squeal_samples[44519]=16231;
squeal_samples[44520]=18564;
squeal_samples[44521]=20786;
squeal_samples[44522]=22923;
squeal_samples[44523]=24956;
squeal_samples[44524]=26898;
squeal_samples[44525]=28758;
squeal_samples[44526]=30527;
squeal_samples[44527]=32225;
squeal_samples[44528]=33843;
squeal_samples[44529]=35386;
squeal_samples[44530]=36868;
squeal_samples[44531]=38271;
squeal_samples[44532]=39624;
squeal_samples[44533]=40908;
squeal_samples[44534]=42134;
squeal_samples[44535]=43308;
squeal_samples[44536]=44424;
squeal_samples[44537]=45494;
squeal_samples[44538]=46518;
squeal_samples[44539]=47491;
squeal_samples[44540]=48422;
squeal_samples[44541]=49317;
squeal_samples[44542]=50158;
squeal_samples[44543]=50973;
squeal_samples[44544]=51746;
squeal_samples[44545]=52487;
squeal_samples[44546]=53194;
squeal_samples[44547]=53869;
squeal_samples[44548]=54519;
squeal_samples[44549]=54922;
squeal_samples[44550]=50637;
squeal_samples[44551]=44774;
squeal_samples[44552]=39272;
squeal_samples[44553]=34133;
squeal_samples[44554]=29315;
squeal_samples[44555]=24809;
squeal_samples[44556]=20589;
squeal_samples[44557]=16644;
squeal_samples[44558]=12948;
squeal_samples[44559]=9492;
squeal_samples[44560]=6251;
squeal_samples[44561]=3409;
squeal_samples[44562]=4699;
squeal_samples[44563]=7538;
squeal_samples[44564]=10248;
squeal_samples[44565]=12846;
squeal_samples[44566]=15321;
squeal_samples[44567]=17690;
squeal_samples[44568]=19959;
squeal_samples[44569]=22123;
squeal_samples[44570]=24194;
squeal_samples[44571]=26173;
squeal_samples[44572]=28061;
squeal_samples[44573]=29866;
squeal_samples[44574]=31585;
squeal_samples[44575]=33237;
squeal_samples[44576]=34804;
squeal_samples[44577]=36311;
squeal_samples[44578]=37740;
squeal_samples[44579]=39115;
squeal_samples[44580]=40421;
squeal_samples[44581]=41671;
squeal_samples[44582]=42861;
squeal_samples[44583]=44005;
squeal_samples[44584]=45090;
squeal_samples[44585]=46131;
squeal_samples[44586]=47123;
squeal_samples[44587]=48064;
squeal_samples[44588]=48977;
squeal_samples[44589]=49833;
squeal_samples[44590]=50665;
squeal_samples[44591]=51448;
squeal_samples[44592]=52206;
squeal_samples[44593]=52921;
squeal_samples[44594]=53612;
squeal_samples[44595]=54267;
squeal_samples[44596]=54900;
squeal_samples[44597]=52878;
squeal_samples[44598]=46920;
squeal_samples[44599]=41283;
squeal_samples[44600]=36014;
squeal_samples[44601]=31074;
squeal_samples[44602]=26456;
squeal_samples[44603]=22128;
squeal_samples[44604]=18075;
squeal_samples[44605]=14301;
squeal_samples[44606]=10748;
squeal_samples[44607]=7435;
squeal_samples[44608]=4328;
squeal_samples[44609]=3639;
squeal_samples[44610]=6479;
squeal_samples[44611]=9234;
squeal_samples[44612]=11874;
squeal_samples[44613]=14394;
squeal_samples[44614]=16812;
squeal_samples[44615]=19107;
squeal_samples[44616]=21313;
squeal_samples[44617]=23415;
squeal_samples[44618]=25434;
squeal_samples[44619]=27348;
squeal_samples[44620]=29191;
squeal_samples[44621]=30936;
squeal_samples[44622]=32617;
squeal_samples[44623]=34217;
squeal_samples[44624]=35744;
squeal_samples[44625]=37209;
squeal_samples[44626]=38596;
squeal_samples[44627]=39933;
squeal_samples[44628]=41196;
squeal_samples[44629]=42415;
squeal_samples[44630]=43575;
squeal_samples[44631]=44682;
squeal_samples[44632]=45733;
squeal_samples[44633]=46747;
squeal_samples[44634]=47706;
squeal_samples[44635]=48630;
squeal_samples[44636]=49504;
squeal_samples[44637]=50350;
squeal_samples[44638]=51152;
squeal_samples[44639]=51918;
squeal_samples[44640]=52647;
squeal_samples[44641]=53349;
squeal_samples[44642]=54013;
squeal_samples[44643]=54654;
squeal_samples[44644]=54408;
squeal_samples[44645]=49119;
squeal_samples[44646]=43346;
squeal_samples[44647]=37935;
squeal_samples[44648]=32880;
squeal_samples[44649]=28140;
squeal_samples[44650]=23703;
squeal_samples[44651]=19554;
squeal_samples[44652]=15681;
squeal_samples[44653]=12043;
squeal_samples[44654]=8642;
squeal_samples[44655]=5459;
squeal_samples[44656]=3211;
squeal_samples[44657]=5398;
squeal_samples[44658]=8202;
squeal_samples[44659]=10888;
squeal_samples[44660]=13454;
squeal_samples[44661]=15908;
squeal_samples[44662]=18244;
squeal_samples[44663]=20488;
squeal_samples[44664]=22632;
squeal_samples[44665]=24677;
squeal_samples[44666]=26633;
squeal_samples[44667]=28498;
squeal_samples[44668]=30284;
squeal_samples[44669]=31987;
squeal_samples[44670]=33616;
squeal_samples[44671]=35171;
squeal_samples[44672]=36655;
squeal_samples[44673]=38075;
squeal_samples[44674]=39425;
squeal_samples[44675]=40723;
squeal_samples[44676]=41954;
squeal_samples[44677]=43136;
squeal_samples[44678]=44261;
squeal_samples[44679]=45333;
squeal_samples[44680]=46366;
squeal_samples[44681]=47341;
squeal_samples[44682]=48282;
squeal_samples[44683]=49176;
squeal_samples[44684]=50029;
squeal_samples[44685]=50844;
squeal_samples[44686]=51620;
squeal_samples[44687]=52366;
squeal_samples[44688]=53078;
squeal_samples[44689]=53758;
squeal_samples[44690]=54410;
squeal_samples[44691]=54976;
squeal_samples[44692]=51373;
squeal_samples[44693]=45454;
squeal_samples[44694]=39912;
squeal_samples[44695]=34730;
squeal_samples[44696]=29870;
squeal_samples[44697]=25324;
squeal_samples[44698]=21071;
squeal_samples[44699]=17092;
squeal_samples[44700]=13365;
squeal_samples[44701]=9882;
squeal_samples[44702]=6616;
squeal_samples[44703]=3611;
squeal_samples[44704]=4305;
squeal_samples[44705]=7159;
squeal_samples[44706]=9891;
squeal_samples[44707]=12494;
squeal_samples[44708]=14990;
squeal_samples[44709]=17373;
squeal_samples[44710]=19652;
squeal_samples[44711]=21829;
squeal_samples[44712]=23910;
squeal_samples[44713]=25899;
squeal_samples[44714]=27802;
squeal_samples[44715]=29610;
squeal_samples[44716]=31348;
squeal_samples[44717]=33005;
squeal_samples[44718]=34586;
squeal_samples[44719]=36097;
squeal_samples[44720]=37539;
squeal_samples[44721]=38915;
squeal_samples[44722]=40233;
squeal_samples[44723]=41485;
squeal_samples[44724]=42690;
squeal_samples[44725]=43831;
squeal_samples[44726]=44929;
squeal_samples[44727]=45975;
squeal_samples[44728]=46969;
squeal_samples[44729]=47922;
squeal_samples[44730]=48839;
squeal_samples[44731]=49701;
squeal_samples[44732]=50538;
squeal_samples[44733]=51320;
squeal_samples[44734]=52086;
squeal_samples[44735]=52804;
squeal_samples[44736]=53502;
squeal_samples[44737]=54154;
squeal_samples[44738]=54795;
squeal_samples[44739]=54049;
squeal_samples[44740]=48423;
squeal_samples[44741]=42689;
squeal_samples[44742]=37331;
squeal_samples[44743]=32305;
squeal_samples[44744]=27606;
squeal_samples[44745]=23199;
squeal_samples[44746]=19087;
squeal_samples[44747]=15234;
squeal_samples[44748]=11624;
squeal_samples[44749]=8252;
squeal_samples[44750]=5092;
squeal_samples[44751]=3274;
squeal_samples[44752]=5769;
squeal_samples[44753]=8558;
squeal_samples[44754]=11226;
squeal_samples[44755]=13775;
squeal_samples[44756]=16209;
squeal_samples[44757]=18544;
squeal_samples[44758]=20765;
squeal_samples[44759]=22894;
squeal_samples[44760]=24933;
squeal_samples[44761]=26869;
squeal_samples[44762]=28732;
squeal_samples[44763]=30501;
squeal_samples[44764]=32197;
squeal_samples[44765]=33813;
squeal_samples[44766]=35358;
squeal_samples[44767]=36836;
squeal_samples[44768]=38240;
squeal_samples[44769]=39585;
squeal_samples[44770]=40872;
squeal_samples[44771]=42096;
squeal_samples[44772]=43270;
squeal_samples[44773]=44392;
squeal_samples[44774]=45462;
squeal_samples[44775]=46480;
squeal_samples[44776]=47454;
squeal_samples[44777]=48385;
squeal_samples[44778]=49272;
squeal_samples[44779]=50124;
squeal_samples[44780]=50931;
squeal_samples[44781]=51706;
squeal_samples[44782]=52448;
squeal_samples[44783]=53152;
squeal_samples[44784]=53825;
squeal_samples[44785]=54477;
squeal_samples[44786]=55038;
squeal_samples[44787]=51436;
squeal_samples[44788]=45504;
squeal_samples[44789]=39958;
squeal_samples[44790]=34770;
squeal_samples[44791]=29905;
squeal_samples[44792]=25365;
squeal_samples[44793]=21100;
squeal_samples[44794]=17115;
squeal_samples[44795]=13397;
squeal_samples[44796]=9902;
squeal_samples[44797]=6640;
squeal_samples[44798]=3625;
squeal_samples[44799]=4325;
squeal_samples[44800]=7175;
squeal_samples[44801]=9899;
squeal_samples[44802]=12512;
squeal_samples[44803]=14999;
squeal_samples[44804]=17382;
squeal_samples[44805]=19660;
squeal_samples[44806]=21838;
squeal_samples[44807]=23915;
squeal_samples[44808]=25904;
squeal_samples[44809]=27801;
squeal_samples[44810]=29614;
squeal_samples[44811]=31352;
squeal_samples[44812]=33003;
squeal_samples[44813]=34588;
squeal_samples[44814]=36090;
squeal_samples[44815]=37538;
squeal_samples[44816]=38913;
squeal_samples[44817]=40226;
squeal_samples[44818]=41487;
squeal_samples[44819]=42683;
squeal_samples[44820]=43831;
squeal_samples[44821]=44918;
squeal_samples[44822]=45968;
squeal_samples[44823]=46965;
squeal_samples[44824]=47916;
squeal_samples[44825]=48826;
squeal_samples[44826]=49698;
squeal_samples[44827]=50518;
squeal_samples[44828]=51317;
squeal_samples[44829]=52068;
squeal_samples[44830]=52794;
squeal_samples[44831]=53484;
squeal_samples[44832]=54144;
squeal_samples[44833]=54776;
squeal_samples[44834]=54046;
squeal_samples[44835]=48410;
squeal_samples[44836]=42685;
squeal_samples[44837]=37312;
squeal_samples[44838]=32296;
squeal_samples[44839]=27588;
squeal_samples[44840]=23187;
squeal_samples[44841]=19067;
squeal_samples[44842]=15215;
squeal_samples[44843]=11611;
squeal_samples[44844]=8237;
squeal_samples[44845]=5073;
squeal_samples[44846]=3255;
squeal_samples[44847]=5755;
squeal_samples[44848]=8545;
squeal_samples[44849]=11206;
squeal_samples[44850]=13760;
squeal_samples[44851]=16198;
squeal_samples[44852]=18521;
squeal_samples[44853]=20749;
squeal_samples[44854]=22879;
squeal_samples[44855]=24912;
squeal_samples[44856]=26853;
squeal_samples[44857]=28709;
squeal_samples[44858]=30484;
squeal_samples[44859]=32177;
squeal_samples[44860]=33794;
squeal_samples[44861]=35338;
squeal_samples[44862]=36818;
squeal_samples[44863]=38224;
squeal_samples[44864]=39573;
squeal_samples[44865]=40851;
squeal_samples[44866]=42085;
squeal_samples[44867]=43253;
squeal_samples[44868]=44376;
squeal_samples[44869]=45439;
squeal_samples[44870]=46464;
squeal_samples[44871]=47432;
squeal_samples[44872]=48369;
squeal_samples[44873]=49254;
squeal_samples[44874]=50108;
squeal_samples[44875]=50910;
squeal_samples[44876]=51693;
squeal_samples[44877]=52428;
squeal_samples[44878]=53138;
squeal_samples[44879]=53811;
squeal_samples[44880]=54458;
squeal_samples[44881]=55019;
squeal_samples[44882]=51416;
squeal_samples[44883]=45483;
squeal_samples[44884]=39949;
squeal_samples[44885]=34750;
squeal_samples[44886]=29897;
squeal_samples[44887]=25341;
squeal_samples[44888]=21088;
squeal_samples[44889]=17102;
squeal_samples[44890]=13375;
squeal_samples[44891]=9885;
squeal_samples[44892]=6619;
squeal_samples[44893]=3608;
squeal_samples[44894]=4304;
squeal_samples[44895]=7155;
squeal_samples[44896]=9881;
squeal_samples[44897]=12492;
squeal_samples[44898]=14980;
squeal_samples[44899]=17365;
squeal_samples[44900]=19638;
squeal_samples[44901]=21820;
squeal_samples[44902]=23896;
squeal_samples[44903]=25883;
squeal_samples[44904]=27784;
squeal_samples[44905]=29595;
squeal_samples[44906]=31331;
squeal_samples[44907]=32986;
squeal_samples[44908]=34565;
squeal_samples[44909]=36074;
squeal_samples[44910]=37518;
squeal_samples[44911]=38893;
squeal_samples[44912]=40208;
squeal_samples[44913]=41465;
squeal_samples[44914]=42666;
squeal_samples[44915]=43810;
squeal_samples[44916]=44901;
squeal_samples[44917]=45946;
squeal_samples[44918]=46948;
squeal_samples[44919]=47895;
squeal_samples[44920]=48808;
squeal_samples[44921]=49676;
squeal_samples[44922]=50502;
squeal_samples[44923]=51295;
squeal_samples[44924]=52051;
squeal_samples[44925]=52773;
squeal_samples[44926]=53465;
squeal_samples[44927]=54124;
squeal_samples[44928]=54759;
squeal_samples[44929]=54023;
squeal_samples[44930]=48395;
squeal_samples[44931]=42661;
squeal_samples[44932]=37296;
squeal_samples[44933]=32275;
squeal_samples[44934]=27568;
squeal_samples[44935]=23171;
squeal_samples[44936]=19044;
squeal_samples[44937]=15198;
squeal_samples[44938]=11590;
squeal_samples[44939]=8218;
squeal_samples[44940]=5055;
squeal_samples[44941]=3234;
squeal_samples[44942]=5737;
squeal_samples[44943]=8525;
squeal_samples[44944]=11187;
squeal_samples[44945]=13740;
squeal_samples[44946]=16179;
squeal_samples[44947]=18502;
squeal_samples[44948]=20730;
squeal_samples[44949]=22859;
squeal_samples[44950]=24894;
squeal_samples[44951]=26831;
squeal_samples[44952]=28692;
squeal_samples[44953]=30465;
squeal_samples[44954]=32156;
squeal_samples[44955]=33776;
squeal_samples[44956]=35319;
squeal_samples[44957]=36797;
squeal_samples[44958]=38207;
squeal_samples[44959]=39552;
squeal_samples[44960]=40832;
squeal_samples[44961]=42065;
squeal_samples[44962]=43236;
squeal_samples[44963]=44353;
squeal_samples[44964]=45424;
squeal_samples[44965]=46440;
squeal_samples[44966]=47417;
squeal_samples[44967]=48345;
squeal_samples[44968]=49240;
squeal_samples[44969]=50084;
squeal_samples[44970]=50894;
squeal_samples[44971]=51671;
squeal_samples[44972]=52411;
squeal_samples[44973]=53117;
squeal_samples[44974]=53794;
squeal_samples[44975]=54435;
squeal_samples[44976]=55003;
squeal_samples[44977]=51394;
squeal_samples[44978]=45467;
squeal_samples[44979]=39925;
squeal_samples[44980]=34735;
squeal_samples[44981]=29873;
squeal_samples[44982]=25327;
squeal_samples[44983]=21065;
squeal_samples[44984]=17083;
squeal_samples[44985]=13357;
squeal_samples[44986]=9864;
squeal_samples[44987]=6602;
squeal_samples[44988]=3587;
squeal_samples[44989]=4284;
squeal_samples[44990]=7138;
squeal_samples[44991]=9859;
squeal_samples[44992]=12475;
squeal_samples[44993]=14960;
squeal_samples[44994]=17344;
squeal_samples[44995]=19620;
squeal_samples[44996]=21801;
squeal_samples[44997]=23875;
squeal_samples[44998]=25867;
squeal_samples[44999]=27760;
squeal_samples[45000]=29579;
squeal_samples[45001]=31309;
squeal_samples[45002]=32970;
squeal_samples[45003]=34543;
squeal_samples[45004]=36057;
squeal_samples[45005]=37495;
squeal_samples[45006]=38877;
squeal_samples[45007]=40187;
squeal_samples[45008]=41447;
squeal_samples[45009]=42646;
squeal_samples[45010]=43791;
squeal_samples[45011]=44881;
squeal_samples[45012]=45928;
squeal_samples[45013]=46927;
squeal_samples[45014]=47877;
squeal_samples[45015]=48788;
squeal_samples[45016]=49657;
squeal_samples[45017]=50484;
squeal_samples[45018]=51273;
squeal_samples[45019]=52035;
squeal_samples[45020]=52750;
squeal_samples[45021]=53449;
squeal_samples[45022]=54104;
squeal_samples[45023]=54738;
squeal_samples[45024]=54007;
squeal_samples[45025]=48372;
squeal_samples[45026]=42644;
squeal_samples[45027]=37277;
squeal_samples[45028]=32254;
squeal_samples[45029]=27551;
squeal_samples[45030]=23150;
squeal_samples[45031]=19025;
squeal_samples[45032]=15179;
squeal_samples[45033]=11571;
squeal_samples[45034]=8198;
squeal_samples[45035]=5037;
squeal_samples[45036]=3214;
squeal_samples[45037]=5717;
squeal_samples[45038]=8506;
squeal_samples[45039]=11168;
squeal_samples[45040]=13721;
squeal_samples[45041]=16160;
squeal_samples[45042]=18482;
squeal_samples[45043]=20710;
squeal_samples[45044]=22841;
squeal_samples[45045]=24873;
squeal_samples[45046]=26814;
squeal_samples[45047]=28671;
squeal_samples[45048]=30445;
squeal_samples[45049]=32139;
squeal_samples[45050]=33754;
squeal_samples[45051]=35301;
squeal_samples[45052]=36778;
squeal_samples[45053]=38186;
squeal_samples[45054]=39534;
squeal_samples[45055]=40813;
squeal_samples[45056]=42045;
squeal_samples[45057]=43216;
squeal_samples[45058]=44335;
squeal_samples[45059]=45402;
squeal_samples[45060]=46425;
squeal_samples[45061]=47394;
squeal_samples[45062]=48328;
squeal_samples[45063]=49219;
squeal_samples[45064]=50065;
squeal_samples[45065]=50875;
squeal_samples[45066]=51652;
squeal_samples[45067]=52391;
squeal_samples[45068]=53098;
squeal_samples[45069]=53775;
squeal_samples[45070]=54415;
squeal_samples[45071]=54985;
squeal_samples[45072]=51373;
squeal_samples[45073]=45449;
squeal_samples[45074]=39905;
squeal_samples[45075]=34716;
squeal_samples[45076]=29855;
squeal_samples[45077]=25304;
squeal_samples[45078]=21050;
squeal_samples[45079]=17061;
squeal_samples[45080]=13338;
squeal_samples[45081]=9846;
squeal_samples[45082]=6581;
squeal_samples[45083]=3568;
squeal_samples[45084]=4267;
squeal_samples[45085]=7113;
squeal_samples[45086]=9846;
squeal_samples[45087]=12451;
squeal_samples[45088]=14943;
squeal_samples[45089]=17324;
squeal_samples[45090]=19600;
squeal_samples[45091]=21781;
squeal_samples[45092]=23858;
squeal_samples[45093]=25844;
squeal_samples[45094]=27745;
squeal_samples[45095]=29555;
squeal_samples[45096]=31294;
squeal_samples[45097]=32947;
squeal_samples[45098]=34527;
squeal_samples[45099]=36034;
squeal_samples[45100]=37478;
squeal_samples[45101]=38856;
squeal_samples[45102]=40169;
squeal_samples[45103]=41428;
squeal_samples[45104]=42625;
squeal_samples[45105]=43772;
squeal_samples[45106]=44861;
squeal_samples[45107]=45910;
squeal_samples[45108]=46907;
squeal_samples[45109]=47856;
squeal_samples[45110]=48772;
squeal_samples[45111]=49634;
squeal_samples[45112]=50467;
squeal_samples[45113]=51251;
squeal_samples[45114]=52016;
squeal_samples[45115]=52732;
squeal_samples[45116]=53428;
squeal_samples[45117]=54083;
squeal_samples[45118]=54720;
squeal_samples[45119]=54463;
squeal_samples[45120]=49163;
squeal_samples[45121]=43386;
squeal_samples[45122]=37967;
squeal_samples[45123]=32899;
squeal_samples[45124]=28155;
squeal_samples[45125]=23715;
squeal_samples[45126]=19557;
squeal_samples[45127]=15673;
squeal_samples[45128]=12031;
squeal_samples[45129]=8624;
squeal_samples[45130]=5434;
squeal_samples[45131]=3185;
squeal_samples[45132]=5370;
squeal_samples[45133]=8172;
squeal_samples[45134]=10855;
squeal_samples[45135]=13414;
squeal_samples[45136]=15868;
squeal_samples[45137]=18202;
squeal_samples[45138]=20446;
squeal_samples[45139]=22584;
squeal_samples[45140]=24623;
squeal_samples[45141]=26582;
squeal_samples[45142]=28440;
squeal_samples[45143]=30229;
squeal_samples[45144]=31927;
squeal_samples[45145]=33556;
squeal_samples[45146]=35110;
squeal_samples[45147]=36587;
squeal_samples[45148]=38012;
squeal_samples[45149]=39362;
squeal_samples[45150]=40651;
squeal_samples[45151]=41887;
squeal_samples[45152]=43063;
squeal_samples[45153]=44194;
squeal_samples[45154]=45261;
squeal_samples[45155]=46293;
squeal_samples[45156]=47264;
squeal_samples[45157]=48208;
squeal_samples[45158]=49093;
squeal_samples[45159]=49951;
squeal_samples[45160]=50761;
squeal_samples[45161]=51546;
squeal_samples[45162]=52285;
squeal_samples[45163]=52995;
squeal_samples[45164]=53680;
squeal_samples[45165]=54324;
squeal_samples[45166]=54946;
squeal_samples[45167]=52922;
squeal_samples[45168]=46946;
squeal_samples[45169]=41309;
squeal_samples[45170]=36016;
squeal_samples[45171]=31082;
squeal_samples[45172]=26445;
squeal_samples[45173]=22116;
squeal_samples[45174]=18064;
squeal_samples[45175]=14273;
squeal_samples[45176]=10724;
squeal_samples[45177]=7395;
squeal_samples[45178]=4292;
squeal_samples[45179]=3590;
squeal_samples[45180]=6430;
squeal_samples[45181]=9181;
squeal_samples[45182]=11820;
squeal_samples[45183]=14341;
squeal_samples[45184]=16751;
squeal_samples[45185]=19044;
squeal_samples[45186]=21252;
squeal_samples[45187]=23348;
squeal_samples[45188]=25364;
squeal_samples[45189]=27281;
squeal_samples[45190]=29111;
squeal_samples[45191]=30870;
squeal_samples[45192]=32539;
squeal_samples[45193]=34141;
squeal_samples[45194]=35662;
squeal_samples[45195]=37121;
squeal_samples[45196]=38518;
squeal_samples[45197]=39843;
squeal_samples[45198]=41117;
squeal_samples[45199]=42325;
squeal_samples[45200]=43483;
squeal_samples[45201]=44592;
squeal_samples[45202]=45640;
squeal_samples[45203]=46659;
squeal_samples[45204]=47613;
squeal_samples[45205]=48538;
squeal_samples[45206]=49412;
squeal_samples[45207]=50253;
squeal_samples[45208]=51053;
squeal_samples[45209]=51817;
squeal_samples[45210]=52548;
squeal_samples[45211]=53247;
squeal_samples[45212]=53914;
squeal_samples[45213]=54551;
squeal_samples[45214]=54948;
squeal_samples[45215]=50662;
squeal_samples[45216]=44776;
squeal_samples[45217]=39275;
squeal_samples[45218]=34121;
squeal_samples[45219]=29299;
squeal_samples[45220]=24782;
squeal_samples[45221]=20557;
squeal_samples[45222]=16605;
squeal_samples[45223]=12900;
squeal_samples[45224]=9444;
squeal_samples[45225]=6195;
squeal_samples[45226]=3352;
squeal_samples[45227]=4632;
squeal_samples[45228]=7468;
squeal_samples[45229]=10177;
squeal_samples[45230]=12771;
squeal_samples[45231]=15244;
squeal_samples[45232]=17616;
squeal_samples[45233]=19876;
squeal_samples[45234]=22038;
squeal_samples[45235]=24106;
squeal_samples[45236]=26080;
squeal_samples[45237]=27972;
squeal_samples[45238]=29769;
squeal_samples[45239]=31495;
squeal_samples[45240]=33137;
squeal_samples[45241]=34712;
squeal_samples[45242]=36209;
squeal_samples[45243]=37647;
squeal_samples[45244]=39008;
squeal_samples[45245]=40322;
squeal_samples[45246]=41563;
squeal_samples[45247]=42758;
squeal_samples[45248]=43891;
squeal_samples[45249]=44981;
squeal_samples[45250]=46020;
squeal_samples[45251]=47008;
squeal_samples[45252]=47959;
squeal_samples[45253]=48859;
squeal_samples[45254]=49722;
squeal_samples[45255]=50548;
squeal_samples[45256]=51336;
squeal_samples[45257]=52085;
squeal_samples[45258]=52803;
squeal_samples[45259]=53490;
squeal_samples[45260]=54147;
squeal_samples[45261]=54780;
squeal_samples[45262]=54030;
squeal_samples[45263]=48397;
squeal_samples[45264]=42665;
squeal_samples[45265]=37293;
squeal_samples[45266]=32265;
squeal_samples[45267]=27558;
squeal_samples[45268]=23154;
squeal_samples[45269]=19032;
squeal_samples[45270]=15179;
squeal_samples[45271]=11564;
squeal_samples[45272]=8190;
squeal_samples[45273]=5025;
squeal_samples[45274]=3202;
squeal_samples[45275]=5704;
squeal_samples[45276]=8487;
squeal_samples[45277]=11154;
squeal_samples[45278]=13698;
squeal_samples[45279]=16139;
squeal_samples[45280]=18461;
squeal_samples[45281]=20688;
squeal_samples[45282]=22815;
squeal_samples[45283]=24849;
squeal_samples[45284]=26790;
squeal_samples[45285]=28642;
squeal_samples[45286]=30420;
squeal_samples[45287]=32109;
squeal_samples[45288]=33731;
squeal_samples[45289]=35266;
squeal_samples[45290]=36746;
squeal_samples[45291]=38155;
squeal_samples[45292]=39499;
squeal_samples[45293]=40783;
squeal_samples[45294]=42006;
squeal_samples[45295]=43179;
squeal_samples[45296]=44297;
squeal_samples[45297]=45365;
squeal_samples[45298]=46385;
squeal_samples[45299]=47363;
squeal_samples[45300]=48291;
squeal_samples[45301]=49179;
squeal_samples[45302]=50031;
squeal_samples[45303]=50832;
squeal_samples[45304]=51613;
squeal_samples[45305]=52345;
squeal_samples[45306]=53056;
squeal_samples[45307]=53730;
squeal_samples[45308]=54373;
squeal_samples[45309]=54993;
squeal_samples[45310]=52175;
squeal_samples[45311]=46191;
squeal_samples[45312]=40598;
squeal_samples[45313]=35354;
squeal_samples[45314]=30454;
squeal_samples[45315]=25864;
squeal_samples[45316]=21564;
squeal_samples[45317]=17547;
squeal_samples[45318]=13788;
squeal_samples[45319]=10263;
squeal_samples[45320]=6969;
squeal_samples[45321]=3882;
squeal_samples[45322]=3888;
squeal_samples[45323]=6749;
squeal_samples[45324]=9492;
squeal_samples[45325]=12114;
squeal_samples[45326]=14619;
squeal_samples[45327]=17009;
squeal_samples[45328]=19297;
squeal_samples[45329]=21488;
squeal_samples[45330]=23580;
squeal_samples[45331]=25580;
squeal_samples[45332]=27483;
squeal_samples[45333]=29314;
squeal_samples[45334]=31046;
squeal_samples[45335]=32718;
squeal_samples[45336]=34301;
squeal_samples[45337]=35826;
squeal_samples[45338]=37271;
squeal_samples[45339]=38654;
squeal_samples[45340]=39982;
squeal_samples[45341]=41234;
squeal_samples[45342]=42446;
squeal_samples[45343]=43595;
squeal_samples[45344]=44695;
squeal_samples[45345]=45746;
squeal_samples[45346]=46745;
squeal_samples[45347]=47705;
squeal_samples[45348]=48618;
squeal_samples[45349]=49490;
squeal_samples[45350]=50323;
squeal_samples[45351]=51121;
squeal_samples[45352]=51880;
squeal_samples[45353]=52612;
squeal_samples[45354]=53298;
squeal_samples[45355]=53968;
squeal_samples[45356]=54598;
squeal_samples[45357]=54725;
squeal_samples[45358]=49876;
squeal_samples[45359]=44041;
squeal_samples[45360]=38583;
squeal_samples[45361]=33473;
squeal_samples[45362]=28690;
squeal_samples[45363]=24208;
squeal_samples[45364]=20019;
squeal_samples[45365]=16097;
squeal_samples[45366]=12427;
squeal_samples[45367]=8994;
squeal_samples[45368]=5777;
squeal_samples[45369]=3180;
squeal_samples[45370]=4963;
squeal_samples[45371]=7787;
squeal_samples[45372]=10478;
squeal_samples[45373]=13059;
squeal_samples[45374]=15518;
squeal_samples[45375]=17874;
squeal_samples[45376]=20125;
squeal_samples[45377]=22274;
squeal_samples[45378]=24332;
squeal_samples[45379]=26297;
squeal_samples[45380]=28168;
squeal_samples[45381]=29965;
squeal_samples[45382]=31675;
squeal_samples[45383]=33310;
squeal_samples[45384]=34872;
squeal_samples[45385]=36360;
squeal_samples[45386]=37791;
squeal_samples[45387]=39147;
squeal_samples[45388]=40449;
squeal_samples[45389]=41688;
squeal_samples[45390]=42873;
squeal_samples[45391]=44006;
squeal_samples[45392]=45084;
squeal_samples[45393]=46118;
squeal_samples[45394]=47097;
squeal_samples[45395]=48046;
squeal_samples[45396]=48936;
squeal_samples[45397]=49798;
squeal_samples[45398]=50616;
squeal_samples[45399]=51399;
squeal_samples[45400]=52149;
squeal_samples[45401]=52861;
squeal_samples[45402]=53547;
squeal_samples[45403]=54197;
squeal_samples[45404]=54824;
squeal_samples[45405]=53492;
squeal_samples[45406]=47634;
squeal_samples[45407]=41940;
squeal_samples[45408]=36619;
squeal_samples[45409]=31633;
squeal_samples[45410]=26962;
squeal_samples[45411]=22594;
squeal_samples[45412]=18504;
squeal_samples[45413]=14686;
squeal_samples[45414]=11106;
squeal_samples[45415]=7746;
squeal_samples[45416]=4621;
squeal_samples[45417]=3311;
squeal_samples[45418]=6029;
squeal_samples[45419]=8797;
squeal_samples[45420]=11448;
squeal_samples[45421]=13986;
squeal_samples[45422]=16407;
squeal_samples[45423]=18720;
squeal_samples[45424]=20931;
squeal_samples[45425]=23045;
squeal_samples[45426]=25066;
squeal_samples[45427]=26997;
squeal_samples[45428]=28844;
squeal_samples[45429]=30606;
squeal_samples[45430]=32287;
squeal_samples[45431]=33895;
squeal_samples[45432]=35429;
squeal_samples[45433]=36895;
squeal_samples[45434]=38294;
squeal_samples[45435]=39634;
squeal_samples[45436]=40908;
squeal_samples[45437]=42133;
squeal_samples[45438]=43286;
squeal_samples[45439]=44408;
squeal_samples[45440]=45461;
squeal_samples[45441]=46486;
squeal_samples[45442]=47444;
squeal_samples[45443]=48378;
squeal_samples[45444]=49251;
squeal_samples[45445]=50105;
squeal_samples[45446]=50902;
squeal_samples[45447]=51680;
squeal_samples[45448]=52408;
squeal_samples[45449]=53114;
squeal_samples[45450]=53782;
squeal_samples[45451]=54426;
squeal_samples[45452]=55039;
squeal_samples[45453]=52216;
squeal_samples[45454]=46232;
squeal_samples[45455]=40628;
squeal_samples[45456]=35386;
squeal_samples[45457]=30478;
squeal_samples[45458]=25884;
squeal_samples[45459]=21583;
squeal_samples[45460]=17561;
squeal_samples[45461]=13797;
squeal_samples[45462]=10273;
squeal_samples[45463]=6976;
squeal_samples[45464]=3887;
squeal_samples[45465]=3889;
squeal_samples[45466]=6754;
squeal_samples[45467]=9496;
squeal_samples[45468]=12110;
squeal_samples[45469]=14620;
squeal_samples[45470]=17002;
squeal_samples[45471]=19299;
squeal_samples[45472]=21484;
squeal_samples[45473]=23573;
squeal_samples[45474]=25573;
squeal_samples[45475]=27474;
squeal_samples[45476]=29302;
squeal_samples[45477]=31039;
squeal_samples[45478]=32704;
squeal_samples[45479]=34289;
squeal_samples[45480]=35812;
squeal_samples[45481]=37258;
squeal_samples[45482]=38643;
squeal_samples[45483]=39961;
squeal_samples[45484]=41224;
squeal_samples[45485]=42430;
squeal_samples[45486]=43579;
squeal_samples[45487]=44675;
squeal_samples[45488]=45729;
squeal_samples[45489]=46726;
squeal_samples[45490]=47686;
squeal_samples[45491]=48599;
squeal_samples[45492]=49474;
squeal_samples[45493]=50301;
squeal_samples[45494]=51106;
squeal_samples[45495]=51859;
squeal_samples[45496]=52587;
squeal_samples[45497]=53283;
squeal_samples[45498]=53940;
squeal_samples[45499]=54582;
squeal_samples[45500]=54970;
squeal_samples[45501]=50678;
squeal_samples[45502]=44791;
squeal_samples[45503]=39279;
squeal_samples[45504]=34124;
squeal_samples[45505]=29294;
squeal_samples[45506]=24777;
squeal_samples[45507]=20550;
squeal_samples[45508]=16592;
squeal_samples[45509]=12894;
squeal_samples[45510]=9420;
squeal_samples[45511]=6177;
squeal_samples[45512]=3325;
squeal_samples[45513]=4607;
squeal_samples[45514]=7441;
squeal_samples[45515]=10154;
squeal_samples[45516]=12741;
squeal_samples[45517]=15223;
squeal_samples[45518]=17581;
squeal_samples[45519]=19846;
squeal_samples[45520]=22008;
squeal_samples[45521]=24073;
squeal_samples[45522]=26045;
squeal_samples[45523]=27934;
squeal_samples[45524]=29733;
squeal_samples[45525]=31457;
squeal_samples[45526]=33097;
squeal_samples[45527]=34668;
squeal_samples[45528]=36169;
squeal_samples[45529]=37602;
squeal_samples[45530]=38969;
squeal_samples[45531]=40277;
squeal_samples[45532]=41518;
squeal_samples[45533]=42714;
squeal_samples[45534]=43850;
squeal_samples[45535]=44938;
squeal_samples[45536]=45972;
squeal_samples[45537]=46962;
squeal_samples[45538]=47911;
squeal_samples[45539]=48810;
squeal_samples[45540]=49677;
squeal_samples[45541]=50497;
squeal_samples[45542]=51286;
squeal_samples[45543]=52035;
squeal_samples[45544]=52757;
squeal_samples[45545]=53442;
squeal_samples[45546]=54093;
squeal_samples[45547]=54727;
squeal_samples[45548]=54458;
squeal_samples[45549]=49162;
squeal_samples[45550]=43370;
squeal_samples[45551]=37953;
squeal_samples[45552]=32880;
squeal_samples[45553]=28128;
squeal_samples[45554]=23682;
squeal_samples[45555]=19524;
squeal_samples[45556]=15632;
squeal_samples[45557]=11995;
squeal_samples[45558]=8578;
squeal_samples[45559]=5391;
squeal_samples[45560]=3135;
squeal_samples[45561]=5321;
squeal_samples[45562]=8122;
squeal_samples[45563]=10801;
squeal_samples[45564]=13362;
squeal_samples[45565]=15816;
squeal_samples[45566]=18146;
squeal_samples[45567]=20386;
squeal_samples[45568]=22522;
squeal_samples[45569]=24566;
squeal_samples[45570]=26516;
squeal_samples[45571]=28381;
squeal_samples[45572]=30163;
squeal_samples[45573]=31863;
squeal_samples[45574]=33493;
squeal_samples[45575]=35039;
squeal_samples[45576]=36526;
squeal_samples[45577]=37938;
squeal_samples[45578]=39290;
squeal_samples[45579]=40584;
squeal_samples[45580]=41809;
squeal_samples[45581]=42995;
squeal_samples[45582]=44114;
squeal_samples[45583]=45192;
squeal_samples[45584]=46210;
squeal_samples[45585]=47197;
squeal_samples[45586]=48128;
squeal_samples[45587]=49019;
squeal_samples[45588]=49872;
squeal_samples[45589]=50686;
squeal_samples[45590]=51469;
squeal_samples[45591]=52206;
squeal_samples[45592]=52921;
squeal_samples[45593]=53594;
squeal_samples[45594]=54246;
squeal_samples[45595]=54865;
squeal_samples[45596]=53531;
squeal_samples[45597]=47663;
squeal_samples[45598]=41974;
squeal_samples[45599]=36643;
squeal_samples[45600]=31655;
squeal_samples[45601]=26977;
squeal_samples[45602]=22610;
squeal_samples[45603]=18512;
squeal_samples[45604]=14694;
squeal_samples[45605]=11104;
squeal_samples[45606]=7759;
squeal_samples[45607]=4611;
squeal_samples[45608]=3313;
squeal_samples[45609]=6022;
squeal_samples[45610]=8793;
squeal_samples[45611]=11441;
squeal_samples[45612]=13975;
squeal_samples[45613]=16395;
squeal_samples[45614]=18708;
squeal_samples[45615]=20918;
squeal_samples[45616]=23035;
squeal_samples[45617]=25054;
squeal_samples[45618]=26980;
squeal_samples[45619]=28826;
squeal_samples[45620]=30583;
squeal_samples[45621]=32266;
squeal_samples[45622]=33876;
squeal_samples[45623]=35409;
squeal_samples[45624]=36869;
squeal_samples[45625]=38275;
squeal_samples[45626]=39608;
squeal_samples[45627]=40889;
squeal_samples[45628]=42106;
squeal_samples[45629]=43268;
squeal_samples[45630]=44382;
squeal_samples[45631]=45436;
squeal_samples[45632]=46455;
squeal_samples[45633]=47423;
squeal_samples[45634]=48348;
squeal_samples[45635]=49227;
squeal_samples[45636]=50072;
squeal_samples[45637]=50879;
squeal_samples[45638]=51642;
squeal_samples[45639]=52378;
squeal_samples[45640]=53079;
squeal_samples[45641]=53753;
squeal_samples[45642]=54395;
squeal_samples[45643]=55003;
squeal_samples[45644]=52185;
squeal_samples[45645]=46197;
squeal_samples[45646]=40601;
squeal_samples[45647]=35352;
squeal_samples[45648]=30445;
squeal_samples[45649]=25849;
squeal_samples[45650]=21553;
squeal_samples[45651]=17524;
squeal_samples[45652]=13767;
squeal_samples[45653]=10237;
squeal_samples[45654]=6942;
squeal_samples[45655]=3856;
squeal_samples[45656]=3848;
squeal_samples[45657]=6718;
squeal_samples[45658]=9454;
squeal_samples[45659]=12074;
squeal_samples[45660]=14583;
squeal_samples[45661]=16972;
squeal_samples[45662]=19259;
squeal_samples[45663]=21444;
squeal_samples[45664]=23537;
squeal_samples[45665]=25531;
squeal_samples[45666]=27443;
squeal_samples[45667]=29262;
squeal_samples[45668]=31001;
squeal_samples[45669]=32669;
squeal_samples[45670]=34252;
squeal_samples[45671]=35772;
squeal_samples[45672]=37220;
squeal_samples[45673]=38604;
squeal_samples[45674]=39922;
squeal_samples[45675]=41185;
squeal_samples[45676]=42393;
squeal_samples[45677]=43537;
squeal_samples[45678]=44645;
squeal_samples[45679]=45688;
squeal_samples[45680]=46692;
squeal_samples[45681]=47650;
squeal_samples[45682]=48559;
squeal_samples[45683]=49435;
squeal_samples[45684]=50264;
squeal_samples[45685]=51063;
squeal_samples[45686]=51824;
squeal_samples[45687]=52547;
squeal_samples[45688]=53245;
squeal_samples[45689]=53901;
squeal_samples[45690]=54542;
squeal_samples[45691]=54933;
squeal_samples[45692]=50637;
squeal_samples[45693]=44760;
squeal_samples[45694]=39238;
squeal_samples[45695]=34093;
squeal_samples[45696]=29254;
squeal_samples[45697]=24739;
squeal_samples[45698]=20510;
squeal_samples[45699]=16554;
squeal_samples[45700]=12856;
squeal_samples[45701]=9380;
squeal_samples[45702]=6141;
squeal_samples[45703]=3282;
squeal_samples[45704]=4572;
squeal_samples[45705]=7400;
squeal_samples[45706]=10116;
squeal_samples[45707]=12703;
squeal_samples[45708]=15184;
squeal_samples[45709]=17541;
squeal_samples[45710]=19810;
squeal_samples[45711]=21965;
squeal_samples[45712]=24037;
squeal_samples[45713]=26013;
squeal_samples[45714]=27892;
squeal_samples[45715]=29699;
squeal_samples[45716]=31412;
squeal_samples[45717]=33063;
squeal_samples[45718]=34632;
squeal_samples[45719]=36132;
squeal_samples[45720]=37563;
squeal_samples[45721]=38930;
squeal_samples[45722]=40237;
squeal_samples[45723]=41482;
squeal_samples[45724]=42672;
squeal_samples[45725]=43814;
squeal_samples[45726]=44898;
squeal_samples[45727]=45935;
squeal_samples[45728]=46921;
squeal_samples[45729]=47873;
squeal_samples[45730]=48772;
squeal_samples[45731]=49636;
squeal_samples[45732]=50463;
squeal_samples[45733]=51242;
squeal_samples[45734]=52000;
squeal_samples[45735]=52717;
squeal_samples[45736]=53401;
squeal_samples[45737]=54058;
squeal_samples[45738]=54685;
squeal_samples[45739]=54423;
squeal_samples[45740]=49120;
squeal_samples[45741]=43333;
squeal_samples[45742]=37913;
squeal_samples[45743]=32843;
squeal_samples[45744]=28088;
squeal_samples[45745]=23644;
squeal_samples[45746]=19484;
squeal_samples[45747]=15597;
squeal_samples[45748]=11951;
squeal_samples[45749]=8544;
squeal_samples[45750]=5348;
squeal_samples[45751]=3100;
squeal_samples[45752]=5280;
squeal_samples[45753]=8085;
squeal_samples[45754]=10759;
squeal_samples[45755]=13328;
squeal_samples[45756]=15771;
squeal_samples[45757]=18114;
squeal_samples[45758]=20342;
squeal_samples[45759]=22487;
squeal_samples[45760]=24524;
squeal_samples[45761]=26479;
squeal_samples[45762]=28341;
squeal_samples[45763]=30127;
squeal_samples[45764]=31823;
squeal_samples[45765]=33453;
squeal_samples[45766]=35001;
squeal_samples[45767]=36487;
squeal_samples[45768]=37899;
squeal_samples[45769]=39254;
squeal_samples[45770]=40541;
squeal_samples[45771]=41774;
squeal_samples[45772]=42952;
squeal_samples[45773]=44079;
squeal_samples[45774]=45150;
squeal_samples[45775]=46174;
squeal_samples[45776]=47157;
squeal_samples[45777]=48089;
squeal_samples[45778]=48981;
squeal_samples[45779]=49831;
squeal_samples[45780]=50650;
squeal_samples[45781]=51427;
squeal_samples[45782]=52170;
squeal_samples[45783]=52881;
squeal_samples[45784]=53554;
squeal_samples[45785]=54208;
squeal_samples[45786]=54824;
squeal_samples[45787]=54080;
squeal_samples[45788]=48434;
squeal_samples[45789]=42689;
squeal_samples[45790]=37312;
squeal_samples[45791]=32271;
squeal_samples[45792]=27560;
squeal_samples[45793]=23149;
squeal_samples[45794]=19019;
squeal_samples[45795]=15163;
squeal_samples[45796]=11546;
squeal_samples[45797]=8162;
squeal_samples[45798]=4996;
squeal_samples[45799]=3165;
squeal_samples[45800]=5662;
squeal_samples[45801]=8441;
squeal_samples[45802]=11105;
squeal_samples[45803]=13654;
squeal_samples[45804]=16083;
squeal_samples[45805]=18410;
squeal_samples[45806]=20636;
squeal_samples[45807]=22755;
squeal_samples[45808]=24790;
squeal_samples[45809]=26727;
squeal_samples[45810]=28582;
squeal_samples[45811]=30350;
squeal_samples[45812]=32040;
squeal_samples[45813]=33657;
squeal_samples[45814]=35197;
squeal_samples[45815]=36673;
squeal_samples[45816]=38073;
squeal_samples[45817]=39422;
squeal_samples[45818]=40707;
squeal_samples[45819]=41926;
squeal_samples[45820]=43101;
squeal_samples[45821]=44216;
squeal_samples[45822]=45285;
squeal_samples[45823]=46301;
squeal_samples[45824]=47277;
squeal_samples[45825]=48204;
squeal_samples[45826]=49093;
squeal_samples[45827]=49934;
squeal_samples[45828]=50748;
squeal_samples[45829]=51522;
squeal_samples[45830]=52256;
squeal_samples[45831]=52965;
squeal_samples[45832]=53638;
squeal_samples[45833]=54283;
squeal_samples[45834]=54900;
squeal_samples[45835]=53562;
squeal_samples[45836]=47693;
squeal_samples[45837]=41993;
squeal_samples[45838]=36657;
squeal_samples[45839]=31664;
squeal_samples[45840]=26991;
squeal_samples[45841]=22613;
squeal_samples[45842]=18515;
squeal_samples[45843]=14691;
squeal_samples[45844]=11104;
squeal_samples[45845]=7743;
squeal_samples[45846]=4606;
squeal_samples[45847]=3298;
squeal_samples[45848]=6009;
squeal_samples[45849]=8777;
squeal_samples[45850]=11419;
squeal_samples[45851]=13960;
squeal_samples[45852]=16371;
squeal_samples[45853]=18691;
squeal_samples[45854]=20894;
squeal_samples[45855]=23010;
squeal_samples[45856]=25026;
squeal_samples[45857]=26952;
squeal_samples[45858]=28802;
squeal_samples[45859]=30554;
squeal_samples[45860]=32241;
squeal_samples[45861]=33843;
squeal_samples[45862]=35381;
squeal_samples[45863]=36845;
squeal_samples[45864]=38239;
squeal_samples[45865]=39580;
squeal_samples[45866]=40854;
squeal_samples[45867]=42069;
squeal_samples[45868]=43238;
squeal_samples[45869]=44339;
squeal_samples[45870]=45410;
squeal_samples[45871]=46413;
squeal_samples[45872]=47389;
squeal_samples[45873]=48308;
squeal_samples[45874]=49190;
squeal_samples[45875]=50028;
squeal_samples[45876]=50843;
squeal_samples[45877]=51603;
squeal_samples[45878]=52341;
squeal_samples[45879]=53040;
squeal_samples[45880]=53712;
squeal_samples[45881]=54354;
squeal_samples[45882]=54968;
squeal_samples[45883]=52932;
squeal_samples[45884]=46950;
squeal_samples[45885]=41295;
squeal_samples[45886]=36005;
squeal_samples[45887]=31053;
squeal_samples[45888]=26416;
squeal_samples[45889]=22077;
squeal_samples[45890]=18017;
squeal_samples[45891]=14220;
squeal_samples[45892]=10663;
squeal_samples[45893]=7335;
squeal_samples[45894]=4218;
squeal_samples[45895]=3519;
squeal_samples[45896]=6352;
squeal_samples[45897]=9104;
squeal_samples[45898]=11735;
squeal_samples[45899]=14260;
squeal_samples[45900]=16655;
squeal_samples[45901]=18957;
squeal_samples[45902]=21151;
squeal_samples[45903]=23262;
squeal_samples[45904]=25258;
squeal_samples[45905]=27185;
squeal_samples[45906]=29011;
squeal_samples[45907]=30763;
squeal_samples[45908]=32437;
squeal_samples[45909]=34031;
squeal_samples[45910]=35552;
squeal_samples[45911]=37014;
squeal_samples[45912]=38398;
squeal_samples[45913]=39737;
squeal_samples[45914]=40993;
squeal_samples[45915]=42209;
squeal_samples[45916]=43366;
squeal_samples[45917]=44470;
squeal_samples[45918]=45526;
squeal_samples[45919]=46530;
squeal_samples[45920]=47493;
squeal_samples[45921]=48412;
squeal_samples[45922]=49290;
squeal_samples[45923]=50122;
squeal_samples[45924]=50929;
squeal_samples[45925]=51688;
squeal_samples[45926]=52417;
squeal_samples[45927]=53118;
squeal_samples[45928]=53785;
squeal_samples[45929]=54419;
squeal_samples[45930]=55031;
squeal_samples[45931]=52199;
squeal_samples[45932]=46213;
squeal_samples[45933]=40607;
squeal_samples[45934]=35358;
squeal_samples[45935]=30448;
squeal_samples[45936]=25845;
squeal_samples[45937]=21548;
squeal_samples[45938]=17518;
squeal_samples[45939]=13748;
squeal_samples[45940]=10227;
squeal_samples[45941]=6919;
squeal_samples[45942]=3838;
squeal_samples[45943]=3826;
squeal_samples[45944]=6693;
squeal_samples[45945]=9430;
squeal_samples[45946]=12048;
squeal_samples[45947]=14552;
squeal_samples[45948]=16942;
squeal_samples[45949]=19226;
squeal_samples[45950]=21416;
squeal_samples[45951]=23504;
squeal_samples[45952]=25495;
squeal_samples[45953]=27409;
squeal_samples[45954]=29222;
squeal_samples[45955]=30969;
squeal_samples[45956]=32624;
squeal_samples[45957]=34218;
squeal_samples[45958]=35729;
squeal_samples[45959]=37178;
squeal_samples[45960]=38564;
squeal_samples[45961]=39878;
squeal_samples[45962]=41147;
squeal_samples[45963]=42346;
squeal_samples[45964]=43501;
squeal_samples[45965]=44593;
squeal_samples[45966]=45644;
squeal_samples[45967]=46644;
squeal_samples[45968]=47603;
squeal_samples[45969]=48511;
squeal_samples[45970]=49388;
squeal_samples[45971]=50217;
squeal_samples[45972]=51017;
squeal_samples[45973]=51769;
squeal_samples[45974]=52503;
squeal_samples[45975]=53187;
squeal_samples[45976]=53859;
squeal_samples[45977]=54485;
squeal_samples[45978]=55044;
squeal_samples[45979]=51418;
squeal_samples[45980]=45481;
squeal_samples[45981]=39922;
squeal_samples[45982]=34716;
squeal_samples[45983]=29844;
squeal_samples[45984]=25284;
squeal_samples[45985]=21015;
squeal_samples[45986]=17021;
squeal_samples[45987]=13287;
squeal_samples[45988]=9793;
squeal_samples[45989]=6516;
squeal_samples[45990]=3496;
squeal_samples[45991]=4189;
squeal_samples[45992]=7024;
squeal_samples[45993]=9757;
squeal_samples[45994]=12355;
squeal_samples[45995]=14850;
squeal_samples[45996]=17217;
squeal_samples[45997]=19496;
squeal_samples[45998]=21670;
squeal_samples[45999]=23752;
squeal_samples[46000]=25729;
squeal_samples[46001]=27631;
squeal_samples[46002]=29437;
squeal_samples[46003]=31168;
squeal_samples[46004]=32824;
squeal_samples[46005]=34396;
squeal_samples[46006]=35905;
squeal_samples[46007]=37348;
squeal_samples[46008]=38720;
squeal_samples[46009]=40034;
squeal_samples[46010]=41286;
squeal_samples[46011]=42487;
squeal_samples[46012]=43623;
squeal_samples[46013]=44723;
squeal_samples[46014]=45761;
squeal_samples[46015]=46756;
squeal_samples[46016]=47707;
squeal_samples[46017]=48615;
squeal_samples[46018]=49482;
squeal_samples[46019]=50311;
squeal_samples[46020]=51098;
squeal_samples[46021]=51855;
squeal_samples[46022]=52577;
squeal_samples[46023]=53268;
squeal_samples[46024]=53928;
squeal_samples[46025]=54555;
squeal_samples[46026]=54945;
squeal_samples[46027]=50651;
squeal_samples[46028]=44756;
squeal_samples[46029]=39242;
squeal_samples[46030]=34080;
squeal_samples[46031]=29249;
squeal_samples[46032]=24725;
squeal_samples[46033]=20492;
squeal_samples[46034]=16535;
squeal_samples[46035]=12831;
squeal_samples[46036]=9357;
squeal_samples[46037]=6111;
squeal_samples[46038]=3253;
squeal_samples[46039]=4542;
squeal_samples[46040]=7366;
squeal_samples[46041]=10080;
squeal_samples[46042]=12665;
squeal_samples[46043]=15140;
squeal_samples[46044]=17504;
squeal_samples[46045]=19767;
squeal_samples[46046]=21928;
squeal_samples[46047]=23989;
squeal_samples[46048]=25968;
squeal_samples[46049]=27845;
squeal_samples[46050]=29654;
squeal_samples[46051]=31368;
squeal_samples[46052]=33015;
squeal_samples[46053]=34582;
squeal_samples[46054]=36081;
squeal_samples[46055]=37510;
squeal_samples[46056]=38882;
squeal_samples[46057]=40178;
squeal_samples[46058]=41431;
squeal_samples[46059]=42622;
squeal_samples[46060]=43756;
squeal_samples[46061]=44843;
squeal_samples[46062]=45876;
squeal_samples[46063]=46873;
squeal_samples[46064]=47813;
squeal_samples[46065]=48718;
squeal_samples[46066]=49579;
squeal_samples[46067]=50399;
squeal_samples[46068]=51188;
squeal_samples[46069]=51935;
squeal_samples[46070]=52657;
squeal_samples[46071]=53339;
squeal_samples[46072]=53995;
squeal_samples[46073]=54621;
squeal_samples[46074]=54738;
squeal_samples[46075]=49875;
squeal_samples[46076]=44042;
squeal_samples[46077]=38563;
squeal_samples[46078]=33456;
squeal_samples[46079]=28656;
squeal_samples[46080]=24174;
squeal_samples[46081]=19975;
squeal_samples[46082]=16052;
squeal_samples[46083]=12370;
squeal_samples[46084]=8935;
squeal_samples[46085]=5710;
squeal_samples[46086]=3113;
squeal_samples[46087]=4887;
squeal_samples[46088]=7707;
squeal_samples[46089]=10394;
squeal_samples[46090]=12972;
squeal_samples[46091]=15433;
squeal_samples[46092]=17785;
squeal_samples[46093]=20026;
squeal_samples[46094]=22181;
squeal_samples[46095]=24232;
squeal_samples[46096]=26198;
squeal_samples[46097]=28065;
squeal_samples[46098]=29860;
squeal_samples[46099]=31569;
squeal_samples[46100]=33209;
squeal_samples[46101]=34758;
squeal_samples[46102]=36259;
squeal_samples[46103]=37674;
squeal_samples[46104]=39037;
squeal_samples[46105]=40336;
squeal_samples[46106]=41569;
squeal_samples[46107]=42756;
squeal_samples[46108]=43886;
squeal_samples[46109]=44964;
squeal_samples[46110]=45991;
squeal_samples[46111]=46982;
squeal_samples[46112]=47919;
squeal_samples[46113]=48815;
squeal_samples[46114]=49674;
squeal_samples[46115]=50491;
squeal_samples[46116]=51277;
squeal_samples[46117]=52017;
squeal_samples[46118]=52734;
squeal_samples[46119]=53416;
squeal_samples[46120]=54067;
squeal_samples[46121]=54688;
squeal_samples[46122]=54802;
squeal_samples[46123]=49940;
squeal_samples[46124]=44090;
squeal_samples[46125]=38622;
squeal_samples[46126]=33493;
squeal_samples[46127]=28706;
squeal_samples[46128]=24210;
squeal_samples[46129]=20010;
squeal_samples[46130]=16084;
squeal_samples[46131]=12402;
squeal_samples[46132]=8959;
squeal_samples[46133]=5737;
squeal_samples[46134]=3133;
squeal_samples[46135]=4911;
squeal_samples[46136]=7724;
squeal_samples[46137]=10417;
squeal_samples[46138]=12989;
squeal_samples[46139]=15448;
squeal_samples[46140]=17798;
squeal_samples[46141]=20047;
squeal_samples[46142]=22190;
squeal_samples[46143]=24248;
squeal_samples[46144]=26207;
squeal_samples[46145]=28079;
squeal_samples[46146]=29870;
squeal_samples[46147]=31579;
squeal_samples[46148]=33211;
squeal_samples[46149]=34771;
squeal_samples[46150]=36259;
squeal_samples[46151]=37686;
squeal_samples[46152]=39036;
squeal_samples[46153]=40337;
squeal_samples[46154]=41578;
squeal_samples[46155]=42758;
squeal_samples[46156]=43894;
squeal_samples[46157]=44964;
squeal_samples[46158]=45998;
squeal_samples[46159]=46979;
squeal_samples[46160]=47922;
squeal_samples[46161]=48817;
squeal_samples[46162]=49672;
squeal_samples[46163]=50492;
squeal_samples[46164]=51266;
squeal_samples[46165]=52025;
squeal_samples[46166]=52731;
squeal_samples[46167]=53413;
squeal_samples[46168]=54064;
squeal_samples[46169]=54680;
squeal_samples[46170]=54803;
squeal_samples[46171]=49931;
squeal_samples[46172]=44091;
squeal_samples[46173]=38614;
squeal_samples[46174]=33490;
squeal_samples[46175]=28697;
squeal_samples[46176]=24204;
squeal_samples[46177]=20009;
squeal_samples[46178]=16072;
squeal_samples[46179]=12399;
squeal_samples[46180]=8955;
squeal_samples[46181]=5732;
squeal_samples[46182]=3124;
squeal_samples[46183]=4901;
squeal_samples[46184]=7720;
squeal_samples[46185]=10409;
squeal_samples[46186]=12983;
squeal_samples[46187]=15444;
squeal_samples[46188]=17790;
squeal_samples[46189]=20034;
squeal_samples[46190]=22191;
squeal_samples[46191]=24233;
squeal_samples[46192]=26202;
squeal_samples[46193]=28066;
squeal_samples[46194]=29862;
squeal_samples[46195]=31568;
squeal_samples[46196]=33205;
squeal_samples[46197]=34757;
squeal_samples[46198]=36254;
squeal_samples[46199]=37671;
squeal_samples[46200]=39030;
squeal_samples[46201]=40332;
squeal_samples[46202]=41568;
squeal_samples[46203]=42752;
squeal_samples[46204]=43878;
squeal_samples[46205]=44961;
squeal_samples[46206]=45988;
squeal_samples[46207]=46974;
squeal_samples[46208]=47911;
squeal_samples[46209]=48806;
squeal_samples[46210]=49667;
squeal_samples[46211]=50480;
squeal_samples[46212]=51266;
squeal_samples[46213]=52007;
squeal_samples[46214]=52727;
squeal_samples[46215]=53402;
squeal_samples[46216]=54053;
squeal_samples[46217]=54680;
squeal_samples[46218]=54789;
squeal_samples[46219]=49924;
squeal_samples[46220]=44081;
squeal_samples[46221]=38603;
squeal_samples[46222]=33485;
squeal_samples[46223]=28688;
squeal_samples[46224]=24198;
squeal_samples[46225]=19997;
squeal_samples[46226]=16069;
squeal_samples[46227]=12389;
squeal_samples[46228]=8945;
squeal_samples[46229]=5724;
squeal_samples[46230]=3112;
squeal_samples[46231]=4894;
squeal_samples[46232]=7708;
squeal_samples[46233]=10401;
squeal_samples[46234]=12973;
squeal_samples[46235]=15435;
squeal_samples[46236]=17778;
squeal_samples[46237]=20029;
squeal_samples[46238]=22175;
squeal_samples[46239]=24232;
squeal_samples[46240]=26184;
squeal_samples[46241]=28063;
squeal_samples[46242]=29848;
squeal_samples[46243]=31562;
squeal_samples[46244]=33192;
squeal_samples[46245]=34757;
squeal_samples[46246]=36241;
squeal_samples[46247]=37664;
squeal_samples[46248]=39020;
squeal_samples[46249]=40322;
squeal_samples[46250]=41559;
squeal_samples[46251]=42741;
squeal_samples[46252]=43871;
squeal_samples[46253]=44949;
squeal_samples[46254]=45981;
squeal_samples[46255]=46963;
squeal_samples[46256]=47901;
squeal_samples[46257]=48798;
squeal_samples[46258]=49655;
squeal_samples[46259]=50474;
squeal_samples[46260]=51253;
squeal_samples[46261]=52001;
squeal_samples[46262]=52715;
squeal_samples[46263]=53392;
squeal_samples[46264]=54052;
squeal_samples[46265]=54665;
squeal_samples[46266]=54785;
squeal_samples[46267]=49911;
squeal_samples[46268]=44073;
squeal_samples[46269]=38593;
squeal_samples[46270]=33475;
squeal_samples[46271]=28678;
squeal_samples[46272]=24190;
squeal_samples[46273]=19985;
squeal_samples[46274]=16063;
squeal_samples[46275]=12377;
squeal_samples[46276]=8938;
squeal_samples[46277]=5711;
squeal_samples[46278]=3105;
squeal_samples[46279]=4885;
squeal_samples[46280]=7697;
squeal_samples[46281]=10393;
squeal_samples[46282]=12962;
squeal_samples[46283]=15425;
squeal_samples[46284]=17772;
squeal_samples[46285]=20016;
squeal_samples[46286]=22168;
squeal_samples[46287]=24219;
squeal_samples[46288]=26178;
squeal_samples[46289]=28051;
squeal_samples[46290]=29840;
squeal_samples[46291]=31552;
squeal_samples[46292]=33182;
squeal_samples[46293]=34748;
squeal_samples[46294]=36231;
squeal_samples[46295]=37655;
squeal_samples[46296]=39010;
squeal_samples[46297]=40312;
squeal_samples[46298]=41550;
squeal_samples[46299]=42732;
squeal_samples[46300]=43861;
squeal_samples[46301]=44939;
squeal_samples[46302]=45973;
squeal_samples[46303]=46950;
squeal_samples[46304]=47897;
squeal_samples[46305]=48783;
squeal_samples[46306]=49648;
squeal_samples[46307]=50466;
squeal_samples[46308]=51240;
squeal_samples[46309]=51995;
squeal_samples[46310]=52703;
squeal_samples[46311]=53384;
squeal_samples[46312]=54040;
squeal_samples[46313]=54660;
squeal_samples[46314]=54771;
squeal_samples[46315]=49906;
squeal_samples[46316]=44059;
squeal_samples[46317]=38586;
squeal_samples[46318]=33464;
squeal_samples[46319]=28670;
squeal_samples[46320]=24180;
squeal_samples[46321]=19976;
squeal_samples[46322]=16051;
squeal_samples[46323]=12370;
squeal_samples[46324]=8926;
squeal_samples[46325]=5704;
squeal_samples[46326]=3096;
squeal_samples[46327]=4871;
squeal_samples[46328]=7693;
squeal_samples[46329]=10379;
squeal_samples[46330]=12955;
squeal_samples[46331]=15416;
squeal_samples[46332]=17760;
squeal_samples[46333]=20008;
squeal_samples[46334]=22159;
squeal_samples[46335]=24208;
squeal_samples[46336]=26170;
squeal_samples[46337]=28040;
squeal_samples[46338]=29832;
squeal_samples[46339]=31541;
squeal_samples[46340]=33174;
squeal_samples[46341]=34736;
squeal_samples[46342]=36224;
squeal_samples[46343]=37644;
squeal_samples[46344]=39001;
squeal_samples[46345]=40303;
squeal_samples[46346]=41540;
squeal_samples[46347]=42721;
squeal_samples[46348]=43853;
squeal_samples[46349]=44929;
squeal_samples[46350]=45963;
squeal_samples[46351]=46943;
squeal_samples[46352]=47883;
squeal_samples[46353]=48778;
squeal_samples[46354]=49637;
squeal_samples[46355]=50454;
squeal_samples[46356]=51235;
squeal_samples[46357]=51980;
squeal_samples[46358]=52698;
squeal_samples[46359]=53373;
squeal_samples[46360]=54031;
squeal_samples[46361]=54650;
squeal_samples[46362]=54761;
squeal_samples[46363]=49896;
squeal_samples[46364]=44051;
squeal_samples[46365]=38576;
squeal_samples[46366]=33456;
squeal_samples[46367]=28658;
squeal_samples[46368]=24173;
squeal_samples[46369]=19964;
squeal_samples[46370]=16045;
squeal_samples[46371]=12357;
squeal_samples[46372]=8920;
squeal_samples[46373]=5692;
squeal_samples[46374]=3087;
squeal_samples[46375]=4863;
squeal_samples[46376]=7681;
squeal_samples[46377]=10372;
squeal_samples[46378]=12944;
squeal_samples[46379]=15408;
squeal_samples[46380]=17748;
squeal_samples[46381]=20002;
squeal_samples[46382]=22145;
squeal_samples[46383]=24204;
squeal_samples[46384]=26156;
squeal_samples[46385]=28034;
squeal_samples[46386]=29821;
squeal_samples[46387]=31531;
squeal_samples[46388]=33166;
squeal_samples[46389]=34725;
squeal_samples[46390]=36217;
squeal_samples[46391]=37632;
squeal_samples[46392]=38993;
squeal_samples[46393]=40293;
squeal_samples[46394]=41530;
squeal_samples[46395]=42713;
squeal_samples[46396]=43842;
squeal_samples[46397]=44921;
squeal_samples[46398]=45952;
squeal_samples[46399]=46935;
squeal_samples[46400]=47872;
squeal_samples[46401]=48770;
squeal_samples[46402]=49625;
squeal_samples[46403]=50449;
squeal_samples[46404]=51220;
squeal_samples[46405]=51977;
squeal_samples[46406]=52683;
squeal_samples[46407]=53367;
squeal_samples[46408]=54018;
squeal_samples[46409]=54644;
squeal_samples[46410]=54749;
squeal_samples[46411]=49889;
squeal_samples[46412]=44040;
squeal_samples[46413]=38566;
squeal_samples[46414]=33446;
squeal_samples[46415]=28650;
squeal_samples[46416]=24162;
squeal_samples[46417]=19957;
squeal_samples[46418]=16031;
squeal_samples[46419]=12353;
squeal_samples[46420]=8904;
squeal_samples[46421]=5689;
squeal_samples[46422]=3072;
squeal_samples[46423]=4857;
squeal_samples[46424]=7670;
squeal_samples[46425]=10362;
squeal_samples[46426]=12936;
squeal_samples[46427]=15396;
squeal_samples[46428]=17741;
squeal_samples[46429]=19990;
squeal_samples[46430]=22138;
squeal_samples[46431]=24192;
squeal_samples[46432]=26148;
squeal_samples[46433]=28023;
squeal_samples[46434]=29813;
squeal_samples[46435]=31520;
squeal_samples[46436]=33159;
squeal_samples[46437]=34713;
squeal_samples[46438]=36208;
squeal_samples[46439]=37622;
squeal_samples[46440]=38985;
squeal_samples[46441]=40282;
squeal_samples[46442]=41522;
squeal_samples[46443]=42703;
squeal_samples[46444]=43832;
squeal_samples[46445]=44912;
squeal_samples[46446]=45942;
squeal_samples[46447]=46925;
squeal_samples[46448]=47864;
squeal_samples[46449]=48760;
squeal_samples[46450]=49616;
squeal_samples[46451]=50437;
squeal_samples[46452]=51214;
squeal_samples[46453]=51963;
squeal_samples[46454]=52677;
squeal_samples[46455]=53356;
squeal_samples[46456]=54010;
squeal_samples[46457]=54632;
squeal_samples[46458]=54742;
squeal_samples[46459]=49876;
squeal_samples[46460]=44035;
squeal_samples[46461]=38554;
squeal_samples[46462]=33437;
squeal_samples[46463]=28642;
squeal_samples[46464]=24149;
squeal_samples[46465]=19951;
squeal_samples[46466]=16020;
squeal_samples[46467]=12343;
squeal_samples[46468]=8896;
squeal_samples[46469]=5678;
squeal_samples[46470]=3063;
squeal_samples[46471]=4849;
squeal_samples[46472]=7658;
squeal_samples[46473]=10355;
squeal_samples[46474]=12924;
squeal_samples[46475]=15388;
squeal_samples[46476]=17732;
squeal_samples[46477]=19979;
squeal_samples[46478]=22130;
squeal_samples[46479]=24181;
squeal_samples[46480]=26141;
squeal_samples[46481]=28011;
squeal_samples[46482]=29804;
squeal_samples[46483]=31512;
squeal_samples[46484]=33145;
squeal_samples[46485]=34710;
squeal_samples[46486]=36192;
squeal_samples[46487]=37618;
squeal_samples[46488]=38972;
squeal_samples[46489]=40273;
squeal_samples[46490]=41514;
squeal_samples[46491]=42691;
squeal_samples[46492]=43824;
squeal_samples[46493]=44902;
squeal_samples[46494]=45932;
squeal_samples[46495]=46918;
squeal_samples[46496]=47851;
squeal_samples[46497]=48752;
squeal_samples[46498]=49605;
squeal_samples[46499]=50429;
squeal_samples[46500]=51204;
squeal_samples[46501]=51952;
squeal_samples[46502]=52670;
squeal_samples[46503]=53341;
squeal_samples[46504]=54006;
squeal_samples[46505]=54617;
squeal_samples[46506]=55007;
squeal_samples[46507]=50691;
squeal_samples[46508]=44795;
squeal_samples[46509]=39274;
squeal_samples[46510]=34106;
squeal_samples[46511]=29261;
squeal_samples[46512]=24733;
squeal_samples[46513]=20493;
squeal_samples[46514]=16522;
squeal_samples[46515]=12818;
squeal_samples[46516]=9340;
squeal_samples[46517]=6095;
squeal_samples[46518]=3225;
squeal_samples[46519]=4513;
squeal_samples[46520]=7336;
squeal_samples[46521]=10042;
squeal_samples[46522]=12632;
squeal_samples[46523]=15097;
squeal_samples[46524]=17463;
squeal_samples[46525]=19721;
squeal_samples[46526]=21880;
squeal_samples[46527]=23945;
squeal_samples[46528]=25912;
squeal_samples[46529]=27797;
squeal_samples[46530]=29593;
squeal_samples[46531]=31313;
squeal_samples[46532]=32952;
squeal_samples[46533]=34518;
squeal_samples[46534]=36018;
squeal_samples[46535]=37449;
squeal_samples[46536]=38811;
squeal_samples[46537]=40118;
squeal_samples[46538]=41360;
squeal_samples[46539]=42549;
squeal_samples[46540]=43689;
squeal_samples[46541]=44773;
squeal_samples[46542]=45804;
squeal_samples[46543]=46797;
squeal_samples[46544]=47741;
squeal_samples[46545]=48643;
squeal_samples[46546]=49500;
squeal_samples[46547]=50326;
squeal_samples[46548]=51107;
squeal_samples[46549]=51857;
squeal_samples[46550]=52577;
squeal_samples[46551]=53258;
squeal_samples[46552]=53917;
squeal_samples[46553]=54540;
squeal_samples[46554]=55085;
squeal_samples[46555]=51457;
squeal_samples[46556]=45507;
squeal_samples[46557]=39937;
squeal_samples[46558]=34727;
squeal_samples[46559]=29843;
squeal_samples[46560]=25277;
squeal_samples[46561]=21006;
squeal_samples[46562]=17001;
squeal_samples[46563]=13263;
squeal_samples[46564]=9756;
squeal_samples[46565]=6480;
squeal_samples[46566]=3451;
squeal_samples[46567]=4145;
squeal_samples[46568]=6982;
squeal_samples[46569]=9704;
squeal_samples[46570]=12303;
squeal_samples[46571]=14793;
squeal_samples[46572]=17164;
squeal_samples[46573]=19435;
squeal_samples[46574]=21605;
squeal_samples[46575]=23678;
squeal_samples[46576]=25667;
squeal_samples[46577]=27557;
squeal_samples[46578]=29369;
squeal_samples[46579]=31094;
squeal_samples[46580]=32750;
squeal_samples[46581]=34317;
squeal_samples[46582]=35831;
squeal_samples[46583]=37264;
squeal_samples[46584]=38640;
squeal_samples[46585]=39950;
squeal_samples[46586]=41201;
squeal_samples[46587]=42397;
squeal_samples[46588]=43538;
squeal_samples[46589]=44629;
squeal_samples[46590]=45667;
squeal_samples[46591]=46666;
squeal_samples[46592]=47610;
squeal_samples[46593]=48520;
squeal_samples[46594]=49388;
squeal_samples[46595]=50211;
squeal_samples[46596]=51008;
squeal_samples[46597]=51758;
squeal_samples[46598]=52482;
squeal_samples[46599]=53166;
squeal_samples[46600]=53831;
squeal_samples[46601]=54454;
squeal_samples[46602]=55060;
squeal_samples[46603]=52217;
squeal_samples[46604]=46220;
squeal_samples[46605]=40609;
squeal_samples[46606]=35350;
squeal_samples[46607]=30433;
squeal_samples[46608]=25821;
squeal_samples[46609]=21509;
squeal_samples[46610]=17480;
squeal_samples[46611]=13704;
squeal_samples[46612]=10177;
squeal_samples[46613]=6866;
squeal_samples[46614]=3774;
squeal_samples[46615]=3765;
squeal_samples[46616]=6628;
squeal_samples[46617]=9362;
squeal_samples[46618]=11974;
squeal_samples[46619]=14479;
squeal_samples[46620]=16861;
squeal_samples[46621]=19149;
squeal_samples[46622]=21328;
squeal_samples[46623]=23422;
squeal_samples[46624]=25409;
squeal_samples[46625]=27318;
squeal_samples[46626]=29134;
squeal_samples[46627]=30876;
squeal_samples[46628]=32531;
squeal_samples[46629]=34121;
squeal_samples[46630]=35633;
squeal_samples[46631]=37079;
squeal_samples[46632]=38461;
squeal_samples[46633]=39778;
squeal_samples[46634]=41040;
squeal_samples[46635]=42240;
squeal_samples[46636]=43394;
squeal_samples[46637]=44488;
squeal_samples[46638]=45535;
squeal_samples[46639]=46535;
squeal_samples[46640]=47488;
squeal_samples[46641]=48402;
squeal_samples[46642]=49268;
squeal_samples[46643]=50106;
squeal_samples[46644]=50899;
squeal_samples[46645]=51658;
squeal_samples[46646]=52384;
squeal_samples[46647]=53070;
squeal_samples[46648]=53739;
squeal_samples[46649]=54369;
squeal_samples[46650]=54978;
squeal_samples[46651]=52932;
squeal_samples[46652]=46938;
squeal_samples[46653]=41277;
squeal_samples[46654]=35978;
squeal_samples[46655]=31019;
squeal_samples[46656]=26371;
squeal_samples[46657]=22029;
squeal_samples[46658]=17960;
squeal_samples[46659]=14155;
squeal_samples[46660]=10593;
squeal_samples[46661]=7256;
squeal_samples[46662]=4137;
squeal_samples[46663]=3436;
squeal_samples[46664]=6265;
squeal_samples[46665]=9015;
squeal_samples[46666]=11645;
squeal_samples[46667]=14159;
squeal_samples[46668]=16558;
squeal_samples[46669]=18859;
squeal_samples[46670]=21051;
squeal_samples[46671]=23158;
squeal_samples[46672]=25156;
squeal_samples[46673]=27074;
squeal_samples[46674]=28903;
squeal_samples[46675]=30649;
squeal_samples[46676]=32321;
squeal_samples[46677]=33915;
squeal_samples[46678]=35442;
squeal_samples[46679]=36893;
squeal_samples[46680]=38284;
squeal_samples[46681]=39607;
squeal_samples[46682]=40875;
squeal_samples[46683]=42089;
squeal_samples[46684]=43240;
squeal_samples[46685]=44344;
squeal_samples[46686]=45395;
squeal_samples[46687]=46401;
squeal_samples[46688]=47359;
squeal_samples[46689]=48278;
squeal_samples[46690]=49156;
squeal_samples[46691]=49993;
squeal_samples[46692]=50792;
squeal_samples[46693]=51551;
squeal_samples[46694]=52286;
squeal_samples[46695]=52981;
squeal_samples[46696]=53646;
squeal_samples[46697]=54285;
squeal_samples[46698]=54890;
squeal_samples[46699]=53543;
squeal_samples[46700]=47661;
squeal_samples[46701]=41958;
squeal_samples[46702]=36615;
squeal_samples[46703]=31612;
squeal_samples[46704]=26926;
squeal_samples[46705]=22547;
squeal_samples[46706]=18437;
squeal_samples[46707]=14610;
squeal_samples[46708]=11016;
squeal_samples[46709]=7654;
squeal_samples[46710]=4510;
squeal_samples[46711]=3196;
squeal_samples[46712]=5904;
squeal_samples[46713]=8667;
squeal_samples[46714]=11316;
squeal_samples[46715]=13844;
squeal_samples[46716]=16263;
squeal_samples[46717]=18565;
squeal_samples[46718]=20772;
squeal_samples[46719]=22887;
squeal_samples[46720]=24902;
squeal_samples[46721]=26833;
squeal_samples[46722]=28668;
squeal_samples[46723]=30431;
squeal_samples[46724]=32103;
squeal_samples[46725]=33712;
squeal_samples[46726]=35242;
squeal_samples[46727]=36704;
squeal_samples[46728]=38102;
squeal_samples[46729]=39432;
squeal_samples[46730]=40714;
squeal_samples[46731]=41920;
squeal_samples[46732]=43096;
squeal_samples[46733]=44195;
squeal_samples[46734]=45256;
squeal_samples[46735]=46273;
squeal_samples[46736]=47234;
squeal_samples[46737]=48162;
squeal_samples[46738]=49037;
squeal_samples[46739]=49880;
squeal_samples[46740]=50685;
squeal_samples[46741]=51448;
squeal_samples[46742]=52187;
squeal_samples[46743]=52881;
squeal_samples[46744]=53558;
squeal_samples[46745]=54191;
squeal_samples[46746]=54805;
squeal_samples[46747]=54050;
squeal_samples[46748]=48394;
squeal_samples[46749]=42642;
squeal_samples[46750]=37247;
squeal_samples[46751]=32209;
squeal_samples[46752]=27485;
squeal_samples[46753]=23069;
squeal_samples[46754]=18929;
squeal_samples[46755]=15066;
squeal_samples[46756]=11440;
squeal_samples[46757]=8056;
squeal_samples[46758]=4876;
squeal_samples[46759]=3049;
squeal_samples[46760]=5539;
squeal_samples[46761]=8321;
squeal_samples[46762]=10981;
squeal_samples[46763]=13519;
squeal_samples[46764]=15956;
squeal_samples[46765]=18271;
squeal_samples[46766]=20494;
squeal_samples[46767]=22619;
squeal_samples[46768]=24647;
squeal_samples[46769]=26581;
squeal_samples[46770]=28434;
squeal_samples[46771]=30201;
squeal_samples[46772]=31889;
squeal_samples[46773]=33508;
squeal_samples[46774]=35045;
squeal_samples[46775]=36521;
squeal_samples[46776]=37918;
squeal_samples[46777]=39266;
squeal_samples[46778]=40540;
squeal_samples[46779]=41771;
squeal_samples[46780]=42934;
squeal_samples[46781]=44055;
squeal_samples[46782]=45114;
squeal_samples[46783]=46138;
squeal_samples[46784]=47108;
squeal_samples[46785]=48034;
squeal_samples[46786]=48923;
squeal_samples[46787]=49766;
squeal_samples[46788]=50578;
squeal_samples[46789]=51347;
squeal_samples[46790]=52088;
squeal_samples[46791]=52787;
squeal_samples[46792]=53466;
squeal_samples[46793]=54104;
squeal_samples[46794]=54727;
squeal_samples[46795]=54449;
squeal_samples[46796]=49134;
squeal_samples[46797]=43329;
squeal_samples[46798]=37897;
squeal_samples[46799]=32811;
squeal_samples[46800]=28054;
squeal_samples[46801]=23593;
squeal_samples[46802]=19430;
squeal_samples[46803]=15523;
squeal_samples[46804]=11875;
squeal_samples[46805]=8455;
squeal_samples[46806]=5256;
squeal_samples[46807]=2995;
squeal_samples[46808]=5169;
squeal_samples[46809]=7971;
squeal_samples[46810]=10644;
squeal_samples[46811]=13201;
squeal_samples[46812]=15647;
squeal_samples[46813]=17980;
squeal_samples[46814]=20212;
squeal_samples[46815]=22351;
squeal_samples[46816]=24385;
squeal_samples[46817]=26335;
squeal_samples[46818]=28200;
squeal_samples[46819]=29976;
squeal_samples[46820]=31674;
squeal_samples[46821]=33295;
squeal_samples[46822]=34849;
squeal_samples[46823]=36328;
squeal_samples[46824]=37739;
squeal_samples[46825]=39091;
squeal_samples[46826]=40375;
squeal_samples[46827]=41608;
squeal_samples[46828]=42784;
squeal_samples[46829]=43909;
squeal_samples[46830]=44975;
squeal_samples[46831]=46003;
squeal_samples[46832]=46978;
squeal_samples[46833]=47914;
squeal_samples[46834]=48799;
squeal_samples[46835]=49660;
squeal_samples[46836]=50463;
squeal_samples[46837]=51252;
squeal_samples[46838]=51980;
squeal_samples[46839]=52695;
squeal_samples[46840]=53371;
squeal_samples[46841]=54015;
squeal_samples[46842]=54637;
squeal_samples[46843]=55012;
squeal_samples[46844]=50703;
squeal_samples[46845]=44799;
squeal_samples[46846]=39272;
squeal_samples[46847]=34099;
squeal_samples[46848]=29253;
squeal_samples[46849]=24722;
squeal_samples[46850]=20475;
squeal_samples[46851]=16505;
squeal_samples[46852]=12799;
squeal_samples[46853]=9312;
squeal_samples[46854]=6065;
squeal_samples[46855]=3199;
squeal_samples[46856]=4478;
squeal_samples[46857]=7301;
squeal_samples[46858]=10005;
squeal_samples[46859]=12589;
squeal_samples[46860]=15061;
squeal_samples[46861]=17424;
squeal_samples[46862]=19678;
squeal_samples[46863]=21840;
squeal_samples[46864]=23895;
squeal_samples[46865]=25872;
squeal_samples[46866]=27749;
squeal_samples[46867]=29550;
squeal_samples[46868]=31266;
squeal_samples[46869]=32909;
squeal_samples[46870]=34473;
squeal_samples[46871]=35967;
squeal_samples[46872]=37400;
squeal_samples[46873]=38758;
squeal_samples[46874]=40070;
squeal_samples[46875]=41310;
squeal_samples[46876]=42498;
squeal_samples[46877]=43633;
squeal_samples[46878]=44717;
squeal_samples[46879]=45753;
squeal_samples[46880]=46742;
squeal_samples[46881]=47687;
squeal_samples[46882]=48584;
squeal_samples[46883]=49447;
squeal_samples[46884]=50261;
squeal_samples[46885]=51055;
squeal_samples[46886]=51799;
squeal_samples[46887]=52521;
squeal_samples[46888]=53198;
squeal_samples[46889]=53858;
squeal_samples[46890]=54482;
squeal_samples[46891]=55079;
squeal_samples[46892]=52242;
squeal_samples[46893]=46228;
squeal_samples[46894]=40621;
squeal_samples[46895]=35350;
squeal_samples[46896]=30431;
squeal_samples[46897]=25818;
squeal_samples[46898]=21507;
squeal_samples[46899]=17470;
squeal_samples[46900]=13692;
squeal_samples[46901]=10162;
squeal_samples[46902]=6848;
squeal_samples[46903]=3754;
squeal_samples[46904]=3741;
squeal_samples[46905]=6604;
squeal_samples[46906]=9336;
squeal_samples[46907]=11951;
squeal_samples[46908]=14448;
squeal_samples[46909]=16831;
squeal_samples[46910]=19120;
squeal_samples[46911]=21298;
squeal_samples[46912]=23386;
squeal_samples[46913]=25375;
squeal_samples[46914]=27282;
squeal_samples[46915]=29097;
squeal_samples[46916]=30839;
squeal_samples[46917]=32491;
squeal_samples[46918]=34085;
squeal_samples[46919]=35589;
squeal_samples[46920]=37040;
squeal_samples[46921]=38418;
squeal_samples[46922]=39740;
squeal_samples[46923]=40996;
squeal_samples[46924]=42197;
squeal_samples[46925]=43345;
squeal_samples[46926]=44443;
squeal_samples[46927]=45489;
squeal_samples[46928]=46488;
squeal_samples[46929]=47443;
squeal_samples[46930]=48353;
squeal_samples[46931]=49225;
squeal_samples[46932]=50052;
squeal_samples[46933]=50855;
squeal_samples[46934]=51605;
squeal_samples[46935]=52331;
squeal_samples[46936]=53025;
squeal_samples[46937]=53687;
squeal_samples[46938]=54317;
squeal_samples[46939]=54925;
squeal_samples[46940]=53571;
squeal_samples[46941]=47688;
squeal_samples[46942]=41978;
squeal_samples[46943]=36624;
squeal_samples[46944]=31621;
squeal_samples[46945]=26932;
squeal_samples[46946]=22553;
squeal_samples[46947]=18440;
squeal_samples[46948]=14609;
squeal_samples[46949]=11013;
squeal_samples[46950]=7644;
squeal_samples[46951]=4501;
squeal_samples[46952]=3181;
squeal_samples[46953]=5888;
squeal_samples[46954]=8653;
squeal_samples[46955]=11294;
squeal_samples[46956]=13826;
squeal_samples[46957]=16241;
squeal_samples[46958]=18544;
squeal_samples[46959]=20754;
squeal_samples[46960]=22863;
squeal_samples[46961]=24880;
squeal_samples[46962]=26803;
squeal_samples[46963]=28647;
squeal_samples[46964]=30400;
squeal_samples[46965]=32082;
squeal_samples[46966]=33677;
squeal_samples[46967]=35212;
squeal_samples[46968]=36673;
squeal_samples[46969]=38070;
squeal_samples[46970]=39402;
squeal_samples[46971]=40680;
squeal_samples[46972]=41893;
squeal_samples[46973]=43055;
squeal_samples[46974]=44160;
squeal_samples[46975]=45227;
squeal_samples[46976]=46230;
squeal_samples[46977]=47206;
squeal_samples[46978]=48116;
squeal_samples[46979]=49009;
squeal_samples[46980]=49836;
squeal_samples[46981]=50653;
squeal_samples[46982]=51408;
squeal_samples[46983]=52151;
squeal_samples[46984]=52841;
squeal_samples[46985]=53512;
squeal_samples[46986]=54156;
squeal_samples[46987]=54767;
squeal_samples[46988]=54489;
squeal_samples[46989]=49172;
squeal_samples[46990]=43354;
squeal_samples[46991]=37922;
squeal_samples[46992]=32830;
squeal_samples[46993]=28070;
squeal_samples[46994]=23611;
squeal_samples[46995]=19439;
squeal_samples[46996]=15530;
squeal_samples[46997]=11880;
squeal_samples[46998]=8453;
squeal_samples[46999]=5259;
squeal_samples[47000]=2986;
squeal_samples[47001]=5172;
squeal_samples[47002]=7965;
squeal_samples[47003]=10636;
squeal_samples[47004]=13194;
squeal_samples[47005]=15638;
squeal_samples[47006]=17971;
squeal_samples[47007]=20201;
squeal_samples[47008]=22333;
squeal_samples[47009]=24376;
squeal_samples[47010]=26324;
squeal_samples[47011]=28177;
squeal_samples[47012]=29961;
squeal_samples[47013]=31657;
squeal_samples[47014]=33278;
squeal_samples[47015]=34829;
squeal_samples[47016]=36304;
squeal_samples[47017]=37719;
squeal_samples[47018]=39070;
squeal_samples[47019]=40352;
squeal_samples[47020]=41587;
squeal_samples[47021]=42757;
squeal_samples[47022]=43880;
squeal_samples[47023]=44957;
squeal_samples[47024]=45972;
squeal_samples[47025]=46955;
squeal_samples[47026]=47882;
squeal_samples[47027]=48778;
squeal_samples[47028]=49625;
squeal_samples[47029]=50439;
squeal_samples[47030]=51211;
squeal_samples[47031]=51960;
squeal_samples[47032]=52664;
squeal_samples[47033]=53339;
squeal_samples[47034]=53989;
squeal_samples[47035]=54603;
squeal_samples[47036]=54981;
squeal_samples[47037]=50671;
squeal_samples[47038]=44764;
squeal_samples[47039]=39242;
squeal_samples[47040]=34065;
squeal_samples[47041]=29222;
squeal_samples[47042]=24689;
squeal_samples[47043]=20442;
squeal_samples[47044]=16473;
squeal_samples[47045]=12760;
squeal_samples[47046]=9281;
squeal_samples[47047]=6032;
squeal_samples[47048]=3161;
squeal_samples[47049]=4444;
squeal_samples[47050]=7265;
squeal_samples[47051]=9971;
squeal_samples[47052]=12558;
squeal_samples[47053]=15028;
squeal_samples[47054]=17383;
squeal_samples[47055]=19646;
squeal_samples[47056]=21800;
squeal_samples[47057]=23865;
squeal_samples[47058]=25827;
squeal_samples[47059]=27716;
squeal_samples[47060]=29515;
squeal_samples[47061]=31230;
squeal_samples[47062]=32869;
squeal_samples[47063]=34436;
squeal_samples[47064]=35935;
squeal_samples[47065]=37360;
squeal_samples[47066]=38729;
squeal_samples[47067]=40030;
squeal_samples[47068]=41272;
squeal_samples[47069]=42462;
squeal_samples[47070]=43592;
squeal_samples[47071]=44682;
squeal_samples[47072]=45714;
squeal_samples[47073]=46706;
squeal_samples[47074]=47644;
squeal_samples[47075]=48553;
squeal_samples[47076]=49402;
squeal_samples[47077]=50235;
squeal_samples[47078]=51013;
squeal_samples[47079]=51763;
squeal_samples[47080]=52482;
squeal_samples[47081]=53166;
squeal_samples[47082]=53820;
squeal_samples[47083]=54444;
squeal_samples[47084]=55044;
squeal_samples[47085]=52199;
squeal_samples[47086]=46196;
squeal_samples[47087]=40576;
squeal_samples[47088]=35320;
squeal_samples[47089]=30387;
squeal_samples[47090]=25784;
squeal_samples[47091]=21468;
squeal_samples[47092]=17431;
squeal_samples[47093]=13657;
squeal_samples[47094]=10120;
squeal_samples[47095]=6814;
squeal_samples[47096]=3713;
squeal_samples[47097]=3706;
squeal_samples[47098]=6563;
squeal_samples[47099]=9302;
squeal_samples[47100]=11909;
squeal_samples[47101]=14414;
squeal_samples[47102]=16790;
squeal_samples[47103]=19085;
squeal_samples[47104]=21257;
squeal_samples[47105]=23352;
squeal_samples[47106]=25333;
squeal_samples[47107]=27247;
squeal_samples[47108]=29059;
squeal_samples[47109]=30799;
squeal_samples[47110]=32458;
squeal_samples[47111]=34040;
squeal_samples[47112]=35558;
squeal_samples[47113]=36997;
squeal_samples[47114]=38384;
squeal_samples[47115]=39699;
squeal_samples[47116]=40961;
squeal_samples[47117]=42157;
squeal_samples[47118]=43309;
squeal_samples[47119]=44404;
squeal_samples[47120]=45451;
squeal_samples[47121]=46450;
squeal_samples[47122]=47406;
squeal_samples[47123]=48315;
squeal_samples[47124]=49187;
squeal_samples[47125]=50013;
squeal_samples[47126]=50818;
squeal_samples[47127]=51566;
squeal_samples[47128]=52294;
squeal_samples[47129]=52989;
squeal_samples[47130]=53644;
squeal_samples[47131]=54285;
squeal_samples[47132]=54882;
squeal_samples[47133]=53537;
squeal_samples[47134]=47649;
squeal_samples[47135]=41940;
squeal_samples[47136]=36587;
squeal_samples[47137]=31581;
squeal_samples[47138]=26897;
squeal_samples[47139]=22513;
squeal_samples[47140]=18404;
squeal_samples[47141]=14569;
squeal_samples[47142]=10977;
squeal_samples[47143]=7605;
squeal_samples[47144]=4464;
squeal_samples[47145]=3142;
squeal_samples[47146]=5850;
squeal_samples[47147]=8617;
squeal_samples[47148]=11254;
squeal_samples[47149]=13790;
squeal_samples[47150]=16201;
squeal_samples[47151]=18509;
squeal_samples[47152]=20712;
squeal_samples[47153]=22830;
squeal_samples[47154]=24838;
squeal_samples[47155]=26769;
squeal_samples[47156]=28606;
squeal_samples[47157]=30365;
squeal_samples[47158]=32040;
squeal_samples[47159]=33643;
squeal_samples[47160]=35172;
squeal_samples[47161]=36636;
squeal_samples[47162]=38033;
squeal_samples[47163]=39362;
squeal_samples[47164]=40643;
squeal_samples[47165]=41855;
squeal_samples[47166]=43016;
squeal_samples[47167]=44125;
squeal_samples[47168]=45186;
squeal_samples[47169]=46195;
squeal_samples[47170]=47164;
squeal_samples[47171]=48083;
squeal_samples[47172]=48964;
squeal_samples[47173]=49808;
squeal_samples[47174]=50605;
squeal_samples[47175]=51378;
squeal_samples[47176]=52107;
squeal_samples[47177]=52805;
squeal_samples[47178]=53475;
squeal_samples[47179]=54116;
squeal_samples[47180]=54730;
squeal_samples[47181]=54825;
squeal_samples[47182]=49947;
squeal_samples[47183]=44091;
squeal_samples[47184]=38603;
squeal_samples[47185]=33468;
squeal_samples[47186]=28660;
squeal_samples[47187]=24161;
squeal_samples[47188]=19947;
squeal_samples[47189]=16011;
squeal_samples[47190]=12322;
squeal_samples[47191]=8870;
squeal_samples[47192]=5641;
squeal_samples[47193]=3027;
squeal_samples[47194]=4801;
squeal_samples[47195]=7611;
squeal_samples[47196]=10301;
squeal_samples[47197]=12872;
squeal_samples[47198]=15324;
squeal_samples[47199]=17672;
squeal_samples[47200]=19913;
squeal_samples[47201]=22057;
squeal_samples[47202]=24109;
squeal_samples[47203]=26064;
squeal_samples[47204]=27933;
squeal_samples[47205]=29722;
squeal_samples[47206]=31429;
squeal_samples[47207]=33056;
squeal_samples[47208]=34617;
squeal_samples[47209]=36098;
squeal_samples[47210]=37526;
squeal_samples[47211]=38875;
squeal_samples[47212]=40178;
squeal_samples[47213]=41410;
squeal_samples[47214]=42592;
squeal_samples[47215]=43715;
squeal_samples[47216]=44795;
squeal_samples[47217]=45820;
squeal_samples[47218]=46809;
squeal_samples[47219]=47740;
squeal_samples[47220]=48643;
squeal_samples[47221]=49489;
squeal_samples[47222]=50314;
squeal_samples[47223]=51087;
squeal_samples[47224]=51833;
squeal_samples[47225]=52545;
squeal_samples[47226]=53225;
squeal_samples[47227]=53879;
squeal_samples[47228]=54494;
squeal_samples[47229]=55094;
squeal_samples[47230]=52246;
squeal_samples[47231]=46237;
squeal_samples[47232]=40616;
squeal_samples[47233]=35346;
squeal_samples[47234]=30422;
squeal_samples[47235]=25809;
squeal_samples[47236]=21487;
squeal_samples[47237]=17455;
squeal_samples[47238]=13667;
squeal_samples[47239]=10134;
squeal_samples[47240]=6819;
squeal_samples[47241]=3728;
squeal_samples[47242]=3704;
squeal_samples[47243]=6573;
squeal_samples[47244]=9295;
squeal_samples[47245]=11914;
squeal_samples[47246]=14406;
squeal_samples[47247]=16796;
squeal_samples[47248]=19075;
squeal_samples[47249]=21260;
squeal_samples[47250]=23336;
squeal_samples[47251]=25334;
squeal_samples[47252]=27235;
squeal_samples[47253]=29056;
squeal_samples[47254]=30788;
squeal_samples[47255]=32449;
squeal_samples[47256]=34026;
squeal_samples[47257]=35547;
squeal_samples[47258]=36984;
squeal_samples[47259]=38372;
squeal_samples[47260]=39686;
squeal_samples[47261]=40945;
squeal_samples[47262]=42143;
squeal_samples[47263]=43292;
squeal_samples[47264]=44386;
squeal_samples[47265]=45434;
squeal_samples[47266]=46432;
squeal_samples[47267]=47388;
squeal_samples[47268]=48298;
squeal_samples[47269]=49168;
squeal_samples[47270]=49999;
squeal_samples[47271]=50789;
squeal_samples[47272]=51554;
squeal_samples[47273]=52273;
squeal_samples[47274]=52966;
squeal_samples[47275]=53630;
squeal_samples[47276]=54255;
squeal_samples[47277]=54865;
squeal_samples[47278]=54094;
squeal_samples[47279]=48437;
squeal_samples[47280]=42666;
squeal_samples[47281]=37278;
squeal_samples[47282]=32222;
squeal_samples[47283]=27488;
squeal_samples[47284]=23071;
squeal_samples[47285]=18919;
squeal_samples[47286]=15056;
squeal_samples[47287]=11422;
squeal_samples[47288]=8031;
squeal_samples[47289]=4850;
squeal_samples[47290]=3014;
squeal_samples[47291]=5499;
squeal_samples[47292]=8278;
squeal_samples[47293]=10934;
squeal_samples[47294]=13477;
squeal_samples[47295]=15909;
squeal_samples[47296]=18223;
squeal_samples[47297]=20441;
squeal_samples[47298]=22567;
squeal_samples[47299]=24587;
squeal_samples[47300]=26525;
squeal_samples[47301]=28369;
squeal_samples[47302]=30143;
squeal_samples[47303]=31827;
squeal_samples[47304]=33435;
squeal_samples[47305]=34976;
squeal_samples[47306]=36445;
squeal_samples[47307]=37851;
squeal_samples[47308]=39190;
squeal_samples[47309]=40471;
squeal_samples[47310]=41694;
squeal_samples[47311]=42855;
squeal_samples[47312]=43979;
squeal_samples[47313]=45036;
squeal_samples[47314]=46055;
squeal_samples[47315]=47026;
squeal_samples[47316]=47952;
squeal_samples[47317]=48839;
squeal_samples[47318]=49684;
squeal_samples[47319]=50488;
squeal_samples[47320]=51261;
squeal_samples[47321]=51997;
squeal_samples[47322]=52703;
squeal_samples[47323]=53372;
squeal_samples[47324]=54020;
squeal_samples[47325]=54628;
squeal_samples[47326]=55005;
squeal_samples[47327]=50685;
squeal_samples[47328]=44777;
squeal_samples[47329]=39246;
squeal_samples[47330]=34066;
squeal_samples[47331]=29222;
squeal_samples[47332]=24684;
squeal_samples[47333]=20436;
squeal_samples[47334]=16459;
squeal_samples[47335]=12746;
squeal_samples[47336]=9264;
squeal_samples[47337]=6011;
squeal_samples[47338]=3144;
squeal_samples[47339]=4420;
squeal_samples[47340]=7239;
squeal_samples[47341]=9949;
squeal_samples[47342]=12526;
squeal_samples[47343]=15000;
squeal_samples[47344]=17354;
squeal_samples[47345]=19615;
squeal_samples[47346]=21766;
squeal_samples[47347]=23834;
squeal_samples[47348]=25799;
squeal_samples[47349]=27681;
squeal_samples[47350]=29474;
squeal_samples[47351]=31195;
squeal_samples[47352]=32834;
squeal_samples[47353]=34396;
squeal_samples[47354]=35894;
squeal_samples[47355]=37320;
squeal_samples[47356]=38682;
squeal_samples[47357]=39990;
squeal_samples[47358]=41232;
squeal_samples[47359]=42420;
squeal_samples[47360]=43554;
squeal_samples[47361]=44634;
squeal_samples[47362]=45669;
squeal_samples[47363]=46659;
squeal_samples[47364]=47601;
squeal_samples[47365]=48503;
squeal_samples[47366]=49361;
squeal_samples[47367]=50180;
squeal_samples[47368]=50967;
squeal_samples[47369]=51719;
squeal_samples[47370]=52428;
squeal_samples[47371]=53118;
squeal_samples[47372]=53765;
squeal_samples[47373]=54399;
squeal_samples[47374]=54990;
squeal_samples[47375]=52944;
squeal_samples[47376]=46935;
squeal_samples[47377]=41272;
squeal_samples[47378]=35959;
squeal_samples[47379]=30992;
squeal_samples[47380]=26338;
squeal_samples[47381]=21988;
squeal_samples[47382]=17912;
squeal_samples[47383]=14104;
squeal_samples[47384]=10538;
squeal_samples[47385]=7194;
squeal_samples[47386]=4073;
squeal_samples[47387]=3363;
squeal_samples[47388]=6190;
squeal_samples[47389]=8936;
squeal_samples[47390]=11563;
squeal_samples[47391]=14075;
squeal_samples[47392]=16474;
squeal_samples[47393]=18766;
squeal_samples[47394]=20963;
squeal_samples[47395]=23055;
squeal_samples[47396]=25060;
squeal_samples[47397]=26975;
squeal_samples[47398]=28803;
squeal_samples[47399]=30551;
squeal_samples[47400]=32217;
squeal_samples[47401]=33812;
squeal_samples[47402]=35330;
squeal_samples[47403]=36786;
squeal_samples[47404]=38172;
squeal_samples[47405]=39499;
squeal_samples[47406]=40761;
squeal_samples[47407]=41971;
squeal_samples[47408]=43128;
squeal_samples[47409]=44226;
squeal_samples[47410]=45283;
squeal_samples[47411]=46282;
squeal_samples[47412]=47248;
squeal_samples[47413]=48155;
squeal_samples[47414]=49038;
squeal_samples[47415]=49864;
squeal_samples[47416]=50667;
squeal_samples[47417]=51430;
squeal_samples[47418]=52161;
squeal_samples[47419]=52855;
squeal_samples[47420]=53518;
squeal_samples[47421]=54154;
squeal_samples[47422]=54761;
squeal_samples[47423]=54484;
squeal_samples[47424]=49153;
squeal_samples[47425]=43343;
squeal_samples[47426]=37899;
squeal_samples[47427]=32807;
squeal_samples[47428]=28038;
squeal_samples[47429]=23577;
squeal_samples[47430]=19399;
squeal_samples[47431]=15498;
squeal_samples[47432]=11834;
squeal_samples[47433]=8417;
squeal_samples[47434]=5206;
squeal_samples[47435]=2944;
squeal_samples[47436]=5117;
squeal_samples[47437]=7912;
squeal_samples[47438]=10581;
squeal_samples[47439]=13138;
squeal_samples[47440]=15584;
squeal_samples[47441]=17911;
squeal_samples[47442]=20142;
squeal_samples[47443]=22278;
squeal_samples[47444]=24310;
squeal_samples[47445]=26262;
squeal_samples[47446]=28115;
squeal_samples[47447]=29895;
squeal_samples[47448]=31590;
squeal_samples[47449]=33210;
squeal_samples[47450]=34758;
squeal_samples[47451]=36238;
squeal_samples[47452]=37649;
squeal_samples[47453]=38999;
squeal_samples[47454]=40287;
squeal_samples[47455]=41510;
squeal_samples[47456]=42690;
squeal_samples[47457]=43811;
squeal_samples[47458]=44881;
squeal_samples[47459]=45901;
squeal_samples[47460]=46877;
squeal_samples[47461]=47812;
squeal_samples[47462]=48699;
squeal_samples[47463]=49556;
squeal_samples[47464]=50361;
squeal_samples[47465]=51140;
squeal_samples[47466]=51878;
squeal_samples[47467]=52584;
squeal_samples[47468]=53267;
squeal_samples[47469]=53906;
squeal_samples[47470]=54526;
squeal_samples[47471]=55067;
squeal_samples[47472]=51429;
squeal_samples[47473]=45467;
squeal_samples[47474]=39889;
squeal_samples[47475]=34671;
squeal_samples[47476]=29781;
squeal_samples[47477]=25210;
squeal_samples[47478]=20919;
squeal_samples[47479]=16916;
squeal_samples[47480]=13169;
squeal_samples[47481]=9658;
squeal_samples[47482]=6375;
squeal_samples[47483]=3350;
squeal_samples[47484]=4025;
squeal_samples[47485]=6872;
squeal_samples[47486]=9587;
squeal_samples[47487]=12183;
squeal_samples[47488]=14668;
squeal_samples[47489]=17037;
squeal_samples[47490]=19311;
squeal_samples[47491]=21473;
squeal_samples[47492]=23548;
squeal_samples[47493]=25528;
squeal_samples[47494]=27424;
squeal_samples[47495]=29230;
squeal_samples[47496]=30954;
squeal_samples[47497]=32607;
squeal_samples[47498]=34175;
squeal_samples[47499]=35684;
squeal_samples[47500]=37116;
squeal_samples[47501]=38494;
squeal_samples[47502]=39797;
squeal_samples[47503]=41052;
squeal_samples[47504]=42246;
squeal_samples[47505]=43384;
squeal_samples[47506]=44475;
squeal_samples[47507]=45519;
squeal_samples[47508]=46506;
squeal_samples[47509]=47459;
squeal_samples[47510]=48356;
squeal_samples[47511]=49232;
squeal_samples[47512]=50053;
squeal_samples[47513]=50841;
squeal_samples[47514]=51599;
squeal_samples[47515]=52312;
squeal_samples[47516]=53007;
squeal_samples[47517]=53657;
squeal_samples[47518]=54291;
squeal_samples[47519]=54893;
squeal_samples[47520]=54118;
squeal_samples[47521]=48454;
squeal_samples[47522]=42680;
squeal_samples[47523]=37285;
squeal_samples[47524]=32228;
squeal_samples[47525]=27497;
squeal_samples[47526]=23071;
squeal_samples[47527]=18918;
squeal_samples[47528]=15049;
squeal_samples[47529]=11417;
squeal_samples[47530]=8012;
squeal_samples[47531]=4840;
squeal_samples[47532]=2996;
squeal_samples[47533]=5487;
squeal_samples[47534]=8262;
squeal_samples[47535]=10921;
squeal_samples[47536]=13455;
squeal_samples[47537]=15886;
squeal_samples[47538]=18200;
squeal_samples[47539]=20420;
squeal_samples[47540]=22537;
squeal_samples[47541]=24567;
squeal_samples[47542]=26494;
squeal_samples[47543]=28348;
squeal_samples[47544]=30110;
squeal_samples[47545]=31797;
squeal_samples[47546]=33411;
squeal_samples[47547]=34942;
squeal_samples[47548]=36417;
squeal_samples[47549]=37813;
squeal_samples[47550]=39156;
squeal_samples[47551]=40433;
squeal_samples[47552]=41658;
squeal_samples[47553]=42819;
squeal_samples[47554]=43942;
squeal_samples[47555]=45002;
squeal_samples[47556]=46017;
squeal_samples[47557]=46990;
squeal_samples[47558]=47916;
squeal_samples[47559]=48803;
squeal_samples[47560]=49641;
squeal_samples[47561]=50454;
squeal_samples[47562]=51222;
squeal_samples[47563]=51958;
squeal_samples[47564]=52658;
squeal_samples[47565]=53332;
squeal_samples[47566]=53978;
squeal_samples[47567]=54585;
squeal_samples[47568]=55126;
squeal_samples[47569]=51480;
squeal_samples[47570]=45518;
squeal_samples[47571]=39938;
squeal_samples[47572]=34708;
squeal_samples[47573]=29821;
squeal_samples[47574]=25240;
squeal_samples[47575]=20953;
squeal_samples[47576]=16946;
squeal_samples[47577]=13190;
squeal_samples[47578]=9682;
squeal_samples[47579]=6390;
squeal_samples[47580]=3366;
squeal_samples[47581]=4039;
squeal_samples[47582]=6884;
squeal_samples[47583]=9597;
squeal_samples[47584]=12190;
squeal_samples[47585]=14683;
squeal_samples[47586]=17044;
squeal_samples[47587]=19320;
squeal_samples[47588]=21481;
squeal_samples[47589]=23557;
squeal_samples[47590]=25531;
squeal_samples[47591]=27426;
squeal_samples[47592]=29226;
squeal_samples[47593]=30955;
squeal_samples[47594]=32600;
squeal_samples[47595]=34178;
squeal_samples[47596]=35675;
squeal_samples[47597]=37120;
squeal_samples[47598]=38486;
squeal_samples[47599]=39798;
squeal_samples[47600]=41043;
squeal_samples[47601]=42237;
squeal_samples[47602]=43384;
squeal_samples[47603]=44465;
squeal_samples[47604]=45512;
squeal_samples[47605]=46499;
squeal_samples[47606]=47448;
squeal_samples[47607]=48352;
squeal_samples[47608]=49215;
squeal_samples[47609]=50048;
squeal_samples[47610]=50832;
squeal_samples[47611]=51585;
squeal_samples[47612]=52304;
squeal_samples[47613]=52994;
squeal_samples[47614]=53649;
squeal_samples[47615]=54278;
squeal_samples[47616]=54879;
squeal_samples[47617]=54105;
squeal_samples[47618]=48439;
squeal_samples[47619]=42670;
squeal_samples[47620]=37268;
squeal_samples[47621]=32217;
squeal_samples[47622]=27478;
squeal_samples[47623]=23056;
squeal_samples[47624]=18906;
squeal_samples[47625]=15030;
squeal_samples[47626]=11402;
squeal_samples[47627]=8003;
squeal_samples[47628]=4822;
squeal_samples[47629]=2981;
squeal_samples[47630]=5465;
squeal_samples[47631]=8246;
squeal_samples[47632]=10900;
squeal_samples[47633]=13444;
squeal_samples[47634]=15871;
squeal_samples[47635]=18183;
squeal_samples[47636]=20405;
squeal_samples[47637]=22520;
squeal_samples[47638]=24545;
squeal_samples[47639]=26479;
squeal_samples[47640]=28326;
squeal_samples[47641]=30094;
squeal_samples[47642]=31777;
squeal_samples[47643]=33391;
squeal_samples[47644]=34926;
squeal_samples[47645]=36396;
squeal_samples[47646]=37801;
squeal_samples[47647]=39142;
squeal_samples[47648]=40415;
squeal_samples[47649]=41643;
squeal_samples[47650]=42809;
squeal_samples[47651]=43920;
squeal_samples[47652]=44985;
squeal_samples[47653]=45998;
squeal_samples[47654]=46971;
squeal_samples[47655]=47898;
squeal_samples[47656]=48783;
squeal_samples[47657]=49624;
squeal_samples[47658]=50433;
squeal_samples[47659]=51206;
squeal_samples[47660]=51936;
squeal_samples[47661]=52649;
squeal_samples[47662]=53309;
squeal_samples[47663]=53962;
squeal_samples[47664]=54565;
squeal_samples[47665]=55108;
squeal_samples[47666]=51461;
squeal_samples[47667]=45500;
squeal_samples[47668]=39917;
squeal_samples[47669]=34692;
squeal_samples[47670]=29800;
squeal_samples[47671]=25223;
squeal_samples[47672]=20933;
squeal_samples[47673]=16927;
squeal_samples[47674]=13174;
squeal_samples[47675]=9665;
squeal_samples[47676]=6374;
squeal_samples[47677]=3345;
squeal_samples[47678]=4027;
squeal_samples[47679]=6867;
squeal_samples[47680]=9575;
squeal_samples[47681]=12174;
squeal_samples[47682]=14661;
squeal_samples[47683]=17030;
squeal_samples[47684]=19297;
squeal_samples[47685]=21466;
squeal_samples[47686]=23534;
squeal_samples[47687]=25517;
squeal_samples[47688]=27403;
squeal_samples[47689]=29218;
squeal_samples[47690]=30930;
squeal_samples[47691]=32587;
squeal_samples[47692]=34155;
squeal_samples[47693]=35660;
squeal_samples[47694]=37098;
squeal_samples[47695]=38469;
squeal_samples[47696]=39779;
squeal_samples[47697]=41024;
squeal_samples[47698]=42220;
squeal_samples[47699]=43362;
squeal_samples[47700]=44450;
squeal_samples[47701]=45488;
squeal_samples[47702]=46487;
squeal_samples[47703]=47424;
squeal_samples[47704]=48337;
squeal_samples[47705]=49199;
squeal_samples[47706]=50030;
squeal_samples[47707]=50813;
squeal_samples[47708]=51568;
squeal_samples[47709]=52284;
squeal_samples[47710]=52977;
squeal_samples[47711]=53628;
squeal_samples[47712]=54261;
squeal_samples[47713]=54860;
squeal_samples[47714]=54086;
squeal_samples[47715]=48423;
squeal_samples[47716]=42647;
squeal_samples[47717]=37254;
squeal_samples[47718]=32194;
squeal_samples[47719]=27463;
squeal_samples[47720]=23035;
squeal_samples[47721]=18889;
squeal_samples[47722]=15010;
squeal_samples[47723]=11385;
squeal_samples[47724]=7981;
squeal_samples[47725]=4807;
squeal_samples[47726]=2959;
squeal_samples[47727]=5450;
squeal_samples[47728]=8224;
squeal_samples[47729]=10884;
squeal_samples[47730]=13422;
squeal_samples[47731]=15855;
squeal_samples[47732]=18163;
squeal_samples[47733]=20387;
squeal_samples[47734]=22501;
squeal_samples[47735]=24527;
squeal_samples[47736]=26460;
squeal_samples[47737]=28307;
squeal_samples[47738]=30076;
squeal_samples[47739]=31757;
squeal_samples[47740]=33375;
squeal_samples[47741]=34905;
squeal_samples[47742]=36378;
squeal_samples[47743]=37783;
squeal_samples[47744]=39122;
squeal_samples[47745]=40397;
squeal_samples[47746]=41625;
squeal_samples[47747]=42788;
squeal_samples[47748]=43903;
squeal_samples[47749]=44967;
squeal_samples[47750]=45977;
squeal_samples[47751]=46954;
squeal_samples[47752]=47879;
squeal_samples[47753]=48763;
squeal_samples[47754]=49608;
squeal_samples[47755]=50413;
squeal_samples[47756]=51187;
squeal_samples[47757]=51919;
squeal_samples[47758]=52627;
squeal_samples[47759]=53294;
squeal_samples[47760]=53942;
squeal_samples[47761]=54546;
squeal_samples[47762]=55091;
squeal_samples[47763]=51439;
squeal_samples[47764]=45484;
squeal_samples[47765]=39897;
squeal_samples[47766]=34675;
squeal_samples[47767]=29780;
squeal_samples[47768]=25205;
squeal_samples[47769]=20913;
squeal_samples[47770]=16910;
squeal_samples[47771]=13153;
squeal_samples[47772]=9649;
squeal_samples[47773]=6354;
squeal_samples[47774]=3327;
squeal_samples[47775]=4008;
squeal_samples[47776]=6847;
squeal_samples[47777]=9557;
squeal_samples[47778]=12158;
squeal_samples[47779]=14640;
squeal_samples[47780]=17011;
squeal_samples[47781]=19280;
squeal_samples[47782]=21445;
squeal_samples[47783]=23519;
squeal_samples[47784]=25494;
squeal_samples[47785]=27389;
squeal_samples[47786]=29195;
squeal_samples[47787]=30915;
squeal_samples[47788]=32567;
squeal_samples[47789]=34134;
squeal_samples[47790]=35647;
squeal_samples[47791]=37073;
squeal_samples[47792]=38456;
squeal_samples[47793]=39755;
squeal_samples[47794]=41011;
squeal_samples[47795]=42195;
squeal_samples[47796]=43350;
squeal_samples[47797]=44425;
squeal_samples[47798]=45475;
squeal_samples[47799]=46464;
squeal_samples[47800]=47408;
squeal_samples[47801]=48317;
squeal_samples[47802]=49181;
squeal_samples[47803]=50012;
squeal_samples[47804]=50793;
squeal_samples[47805]=51550;
squeal_samples[47806]=52266;
squeal_samples[47807]=52956;
squeal_samples[47808]=53613;
squeal_samples[47809]=54239;
squeal_samples[47810]=54842;
squeal_samples[47811]=54069;
squeal_samples[47812]=48402;
squeal_samples[47813]=42630;
squeal_samples[47814]=37234;
squeal_samples[47815]=32176;
squeal_samples[47816]=27444;
squeal_samples[47817]=23017;
squeal_samples[47818]=18869;
squeal_samples[47819]=14993;
squeal_samples[47820]=11364;
squeal_samples[47821]=7965;
squeal_samples[47822]=4787;
squeal_samples[47823]=2940;
squeal_samples[47824]=5432;
squeal_samples[47825]=8205;
squeal_samples[47826]=10865;
squeal_samples[47827]=13405;
squeal_samples[47828]=15835;
squeal_samples[47829]=18145;
squeal_samples[47830]=20367;
squeal_samples[47831]=22484;
squeal_samples[47832]=24507;
squeal_samples[47833]=26442;
squeal_samples[47834]=28289;
squeal_samples[47835]=30056;
squeal_samples[47836]=31739;
squeal_samples[47837]=33356;
squeal_samples[47838]=34886;
squeal_samples[47839]=36361;
squeal_samples[47840]=37763;
squeal_samples[47841]=39104;
squeal_samples[47842]=40379;
squeal_samples[47843]=41604;
squeal_samples[47844]=42773;
squeal_samples[47845]=43883;
squeal_samples[47846]=44946;
squeal_samples[47847]=45963;
squeal_samples[47848]=46930;
squeal_samples[47849]=47865;
squeal_samples[47850]=48741;
squeal_samples[47851]=49591;
squeal_samples[47852]=50392;
squeal_samples[47853]=51171;
squeal_samples[47854]=51899;
squeal_samples[47855]=52608;
squeal_samples[47856]=53276;
squeal_samples[47857]=53922;
squeal_samples[47858]=54529;
squeal_samples[47859]=55071;
squeal_samples[47860]=51422;
squeal_samples[47861]=45464;
squeal_samples[47862]=39879;
squeal_samples[47863]=34656;
squeal_samples[47864]=29762;
squeal_samples[47865]=25185;
squeal_samples[47866]=20898;
squeal_samples[47867]=16886;
squeal_samples[47868]=13139;
squeal_samples[47869]=9627;
squeal_samples[47870]=6337;
squeal_samples[47871]=3309;
squeal_samples[47872]=3988;
squeal_samples[47873]=6829;
squeal_samples[47874]=9538;
squeal_samples[47875]=12139;
squeal_samples[47876]=14622;
squeal_samples[47877]=16992;
squeal_samples[47878]=19262;
squeal_samples[47879]=21425;
squeal_samples[47880]=23501;
squeal_samples[47881]=25476;
squeal_samples[47882]=27368;
squeal_samples[47883]=29179;
squeal_samples[47884]=30895;
squeal_samples[47885]=32546;
squeal_samples[47886]=34121;
squeal_samples[47887]=35621;
squeal_samples[47888]=37062;
squeal_samples[47889]=38430;
squeal_samples[47890]=39742;
squeal_samples[47891]=40987;
squeal_samples[47892]=42182;
squeal_samples[47893]=43326;
squeal_samples[47894]=44411;
squeal_samples[47895]=45453;
squeal_samples[47896]=46446;
squeal_samples[47897]=47389;
squeal_samples[47898]=48298;
squeal_samples[47899]=49163;
squeal_samples[47900]=49993;
squeal_samples[47901]=50775;
squeal_samples[47902]=51528;
squeal_samples[47903]=52251;
squeal_samples[47904]=52933;
squeal_samples[47905]=53597;
squeal_samples[47906]=54218;
squeal_samples[47907]=54824;
squeal_samples[47908]=54533;
squeal_samples[47909]=49197;
squeal_samples[47910]=43378;
squeal_samples[47911]=37927;
squeal_samples[47912]=32825;
squeal_samples[47913]=28055;
squeal_samples[47914]=23578;
squeal_samples[47915]=19400;
squeal_samples[47916]=15489;
squeal_samples[47917]=11824;
squeal_samples[47918]=8397;
squeal_samples[47919]=5185;
squeal_samples[47920]=2913;
squeal_samples[47921]=5090;
squeal_samples[47922]=7877;
squeal_samples[47923]=10548;
squeal_samples[47924]=13098;
squeal_samples[47925]=15539;
squeal_samples[47926]=17865;
squeal_samples[47927]=20100;
squeal_samples[47928]=22226;
squeal_samples[47929]=24261;
squeal_samples[47930]=26210;
squeal_samples[47931]=28065;
squeal_samples[47932]=29841;
squeal_samples[47933]=31533;
squeal_samples[47934]=33155;
squeal_samples[47935]=34702;
squeal_samples[47936]=36177;
squeal_samples[47937]=37588;
squeal_samples[47938]=38934;
squeal_samples[47939]=40217;
squeal_samples[47940]=41447;
squeal_samples[47941]=42621;
squeal_samples[47942]=43741;
squeal_samples[47943]=44808;
squeal_samples[47944]=45828;
squeal_samples[47945]=46808;
squeal_samples[47946]=47735;
squeal_samples[47947]=48634;
squeal_samples[47948]=49471;
squeal_samples[47949]=50289;
squeal_samples[47950]=51058;
squeal_samples[47951]=51803;
squeal_samples[47952]=52505;
squeal_samples[47953]=53183;
squeal_samples[47954]=53831;
squeal_samples[47955]=54444;
squeal_samples[47956]=55039;
squeal_samples[47957]=52974;
squeal_samples[47958]=46967;
squeal_samples[47959]=41288;
squeal_samples[47960]=35972;
squeal_samples[47961]=30993;
squeal_samples[47962]=26334;
squeal_samples[47963]=21973;
squeal_samples[47964]=17893;
squeal_samples[47965]=14075;
squeal_samples[47966]=10511;
squeal_samples[47967]=7155;
squeal_samples[47968]=4033;
squeal_samples[47969]=3314;
squeal_samples[47970]=6142;
squeal_samples[47971]=8886;
squeal_samples[47972]=11508;
squeal_samples[47973]=14020;
squeal_samples[47974]=16413;
squeal_samples[47975]=18709;
squeal_samples[47976]=20899;
squeal_samples[47977]=22992;
squeal_samples[47978]=24997;
squeal_samples[47979]=26905;
squeal_samples[47980]=28735;
squeal_samples[47981]=30475;
squeal_samples[47982]=32144;
squeal_samples[47983]=33731;
squeal_samples[47984]=35252;
squeal_samples[47985]=36704;
squeal_samples[47986]=38089;
squeal_samples[47987]=39411;
squeal_samples[47988]=40678;
squeal_samples[47989]=41884;
squeal_samples[47990]=43038;
squeal_samples[47991]=44136;
squeal_samples[47992]=45190;
squeal_samples[47993]=46195;
squeal_samples[47994]=47153;
squeal_samples[47995]=48068;
squeal_samples[47996]=48937;
squeal_samples[47997]=49779;
squeal_samples[47998]=50571;
squeal_samples[47999]=51338;
