library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity prog is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of prog is
	type rom is array(0 to  12287) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"46",X"39",X"90",X"FC",X"20",X"BA",X"58",X"A6",X"28",X"F0",X"FC",X"A9",X"02",X"85",X"02",X"86",
		X"03",X"A9",X"01",X"20",X"81",X"7A",X"20",X"6A",X"7A",X"A9",X"81",X"AA",X"A0",X"00",X"20",X"8E",
		X"7A",X"A9",X"00",X"20",X"63",X"7A",X"E6",X"C6",X"D0",X"06",X"E6",X"D2",X"A5",X"D2",X"C9",X"04",
		X"24",X"CD",X"10",X"06",X"20",X"D9",X"51",X"4C",X"C5",X"53",X"24",X"CE",X"30",X"2D",X"A5",X"C7",
		X"D0",X"29",X"90",X"1C",X"20",X"E8",X"69",X"A2",X"03",X"AD",X"3C",X"03",X"49",X"80",X"8D",X"3C",
		X"03",X"86",X"D2",X"85",X"C6",X"30",X"09",X"24",X"CE",X"30",X"19",X"A9",X"FF",X"8D",X"4B",X"03",
		X"2C",X"3C",X"03",X"10",X"0F",X"20",X"D9",X"51",X"4C",X"9B",X"54",X"90",X"07",X"24",X"CB",X"30",
		X"03",X"20",X"22",X"6A",X"20",X"6A",X"7A",X"A9",X"7F",X"A2",X"30",X"A0",X"00",X"20",X"8E",X"7A",
		X"A9",X"02",X"20",X"63",X"7A",X"24",X"CE",X"30",X"05",X"A2",X"2E",X"20",X"98",X"6C",X"20",X"C8",
		X"57",X"C6",X"C4",X"A5",X"D1",X"C9",X"FF",X"F0",X"02",X"E6",X"D1",X"A9",X"0A",X"8D",X"6C",X"18",
		X"A9",X"00",X"85",X"10",X"20",X"46",X"59",X"20",X"68",X"52",X"A6",X"10",X"BD",X"70",X"02",X"30",
		X"11",X"20",X"4A",X"5D",X"A6",X"10",X"BD",X"70",X"02",X"20",X"5C",X"5C",X"E6",X"10",X"E6",X"10",
		X"D0",X"E8",X"A5",X"C7",X"F0",X"03",X"4C",X"E9",X"51",X"20",X"D9",X"51",X"20",X"E9",X"6A",X"20",
		X"10",X"68",X"49",X"80",X"38",X"E5",X"2A",X"85",X"16",X"10",X"05",X"18",X"49",X"FF",X"69",X"01",
		X"85",X"D0",X"2C",X"4B",X"03",X"30",X"1B",X"C9",X"02",X"A5",X"24",X"F0",X"06",X"A9",X"20",X"25",
		X"3A",X"F0",X"0F",X"90",X"06",X"A2",X"CC",X"A9",X"34",X"D0",X"04",X"A2",X"00",X"A9",X"35",X"20",
		X"5A",X"7A",X"A5",X"14",X"D0",X"44",X"24",X"CE",X"30",X"1C",X"A5",X"03",X"29",X"F8",X"85",X"3C",
		X"A9",X"02",X"85",X"3B",X"A0",X"35",X"A9",X"00",X"51",X"3B",X"88",X"10",X"FB",X"4A",X"8D",X"ED",
		X"02",X"2C",X"4B",X"03",X"30",X"33",X"A9",X"02",X"25",X"C6",X"F0",X"1E",X"A5",X"D0",X"C9",X"16",
		X"90",X"18",X"A2",X"00",X"20",X"98",X"6C",X"A2",X"06",X"A9",X"6B",X"C5",X"D0",X"90",X"08",X"A2",
		X"02",X"24",X"16",X"10",X"02",X"A2",X"04",X"20",X"98",X"6C",X"A5",X"C8",X"F0",X"0B",X"A5",X"C6",
		X"29",X"04",X"D0",X"05",X"A2",X"12",X"20",X"98",X"6C",X"20",X"2E",X"6D",X"A5",X"CD",X"F0",X"31",
		X"A5",X"C7",X"D0",X"2D",X"2C",X"4B",X"03",X"30",X"28",X"A2",X"14",X"20",X"98",X"6C",X"A5",X"0E",
		X"D0",X"16",X"A5",X"EB",X"29",X"03",X"F0",X"10",X"0A",X"69",X"1E",X"AA",X"20",X"98",X"6C",X"A2",
		X"26",X"20",X"98",X"6C",X"A2",X"28",X"D0",X"02",X"A2",X"16",X"24",X"3A",X"50",X"03",X"20",X"98",
		X"6C",X"20",X"74",X"55",X"2C",X"45",X"03",X"30",X"29",X"A9",X"04",X"85",X"18",X"20",X"45",X"60",
		X"20",X"66",X"6C",X"C6",X"18",X"D0",X"F6",X"24",X"CB",X"30",X"05",X"20",X"B5",X"69",X"90",X"03",
		X"20",X"4E",X"5F",X"20",X"18",X"64",X"20",X"7C",X"67",X"20",X"44",X"5E",X"20",X"D0",X"61",X"4C",
		X"00",X"50",X"AD",X"ED",X"02",X"4A",X"05",X"EF",X"D0",X"F5",X"8D",X"45",X"03",X"A5",X"15",X"09",
		X"02",X"85",X"15",X"A9",X"FF",X"85",X"0F",X"D0",X"E6",X"20",X"6A",X"7A",X"A0",X"00",X"A9",X"7F",
		X"AA",X"20",X"8E",X"7A",X"A9",X"02",X"4C",X"63",X"7A",X"A0",X"00",X"8C",X"27",X"18",X"B9",X"F8",
		X"36",X"BE",X"F9",X"36",X"84",X"08",X"20",X"6E",X"7A",X"A4",X"08",X"C8",X"C8",X"C4",X"C7",X"B0",
		X"61",X"C0",X"10",X"90",X"E9",X"A9",X"2C",X"C5",X"C7",X"B0",X"57",X"A5",X"24",X"D0",X"50",X"85",
		X"C7",X"85",X"C5",X"85",X"12",X"85",X"D1",X"A6",X"CD",X"F0",X"07",X"85",X"CE",X"85",X"C8",X"4C",
		X"44",X"53",X"A9",X"30",X"85",X"C4",X"AD",X"2A",X"18",X"85",X"BC",X"85",X"2D",X"AD",X"2A",X"18",
		X"85",X"31",X"AD",X"2A",X"18",X"29",X"3F",X"85",X"2E",X"AD",X"2A",X"18",X"85",X"32",X"A2",X"00",
		X"20",X"D6",X"68",X"B0",X"ED",X"86",X"C8",X"86",X"C9",X"AD",X"2A",X"18",X"85",X"2A",X"24",X"CB",
		X"10",X"06",X"20",X"E8",X"69",X"4C",X"59",X"51",X"A5",X"14",X"D0",X"03",X"20",X"BE",X"69",X"4C",
		X"59",X"51",X"E6",X"C7",X"E6",X"C7",X"D0",X"F7",X"24",X"CE",X"30",X"20",X"A5",X"03",X"29",X"F8",
		X"85",X"3C",X"A9",X"02",X"85",X"3B",X"A0",X"35",X"A9",X"00",X"38",X"F1",X"3B",X"88",X"10",X"FB",
		X"38",X"ED",X"93",X"74",X"8D",X"70",X"03",X"2C",X"4B",X"03",X"30",X"01",X"60",X"AD",X"49",X"03",
		X"30",X"07",X"C9",X"02",X"90",X"03",X"4C",X"1F",X"53",X"A2",X"00",X"BD",X"70",X"02",X"30",X"04",
		X"E8",X"E8",X"D0",X"F7",X"A9",X"F0",X"8D",X"EA",X"02",X"A0",X"00",X"B9",X"F7",X"3F",X"9D",X"70",
		X"02",X"AD",X"46",X"03",X"9D",X"00",X"02",X"A9",X"00",X"9D",X"38",X"02",X"E8",X"C8",X"A5",X"2A",
		X"9D",X"70",X"02",X"AD",X"47",X"03",X"9D",X"00",X"02",X"A9",X"00",X"9D",X"38",X"02",X"E8",X"C8",
		X"AD",X"49",X"03",X"10",X"10",X"C9",X"FD",X"B0",X"0C",X"AD",X"48",X"03",X"C9",X"B0",X"B0",X"05",
		X"C0",X"03",X"4C",X"E7",X"52",X"C0",X"05",X"90",X"C2",X"AD",X"48",X"03",X"AC",X"49",X"03",X"8D",
		X"E4",X"02",X"8C",X"E5",X"02",X"8D",X"E6",X"02",X"8C",X"E7",X"02",X"18",X"69",X"08",X"8D",X"48",
		X"03",X"90",X"01",X"C8",X"8C",X"49",X"03",X"18",X"AC",X"47",X"03",X"AD",X"46",X"03",X"69",X"40",
		X"8D",X"46",X"03",X"90",X"01",X"C8",X"8C",X"47",X"03",X"A9",X"FF",X"9D",X"70",X"02",X"60",X"A9",
		X"FC",X"8D",X"49",X"03",X"A9",X"00",X"8D",X"46",X"03",X"8D",X"48",X"03",X"8D",X"4B",X"03",X"A9",
		X"04",X"8D",X"47",X"03",X"A9",X"03",X"85",X"D2",X"A9",X"00",X"8D",X"3C",X"03",X"85",X"C6",X"60",
		X"70",X"45",X"44",X"52",X"A2",X"00",X"86",X"D2",X"8E",X"3C",X"03",X"BC",X"00",X"03",X"C4",X"B8",
		X"BD",X"01",X"03",X"E5",X"B9",X"90",X"0A",X"E8",X"E8",X"E8",X"E0",X"1E",X"90",X"ED",X"4C",X"59",
		X"51",X"A9",X"00",X"85",X"C6",X"8D",X"42",X"03",X"8E",X"40",X"03",X"85",X"C8",X"85",X"D4",X"85",
		X"DE",X"A9",X"80",X"20",X"85",X"79",X"A5",X"CD",X"09",X"80",X"85",X"CD",X"A2",X"1B",X"EC",X"40",
		X"03",X"F0",X"23",X"BD",X"FD",X"02",X"9D",X"00",X"03",X"BD",X"FE",X"02",X"9D",X"01",X"03",X"BD",
		X"1B",X"03",X"9D",X"1E",X"03",X"BD",X"1C",X"03",X"9D",X"1F",X"03",X"BD",X"1D",X"03",X"9D",X"20",
		X"03",X"CA",X"CA",X"CA",X"10",X"D8",X"A5",X"B8",X"9D",X"00",X"03",X"A5",X"B9",X"9D",X"01",X"03",
		X"A9",X"04",X"8D",X"41",X"03",X"A9",X"16",X"8D",X"3D",X"03",X"A9",X"4C",X"8D",X"3E",X"03",X"8D",
		X"3F",X"03",X"4C",X"59",X"51",X"A5",X"D2",X"C9",X"04",X"B0",X"77",X"A5",X"EF",X"D0",X"0E",X"A6",
		X"BA",X"F0",X"0A",X"85",X"BA",X"A9",X"02",X"85",X"15",X"A9",X"FF",X"85",X"0F",X"20",X"2E",X"6D",
		X"A2",X"1E",X"20",X"98",X"6C",X"A2",X"08",X"20",X"98",X"6C",X"A2",X"0A",X"20",X"98",X"6C",X"A2",
		X"0C",X"20",X"98",X"6C",X"20",X"65",X"54",X"AD",X"28",X"18",X"8D",X"44",X"03",X"4D",X"43",X"03",
		X"2D",X"44",X"03",X"AE",X"44",X"03",X"8E",X"43",X"03",X"29",X"10",X"F0",X"10",X"AE",X"42",X"03",
		X"E0",X"02",X"B0",X"2E",X"E8",X"8E",X"42",X"03",X"A9",X"16",X"9D",X"3D",X"03",X"20",X"6A",X"7A",
		X"A0",X"00",X"84",X"00",X"A9",X"EE",X"A2",X"EE",X"20",X"8E",X"7A",X"A2",X"00",X"86",X"08",X"BD",
		X"3D",X"03",X"20",X"6A",X"55",X"A6",X"08",X"E8",X"E0",X"03",X"90",X"F1",X"20",X"74",X"55",X"4C",
		X"00",X"50",X"AE",X"40",X"03",X"A0",X"00",X"B9",X"3D",X"03",X"9D",X"1E",X"03",X"C0",X"02",X"90",
		X"10",X"A9",X"03",X"85",X"D2",X"85",X"CD",X"A9",X"81",X"8D",X"3C",X"03",X"85",X"C6",X"4C",X"00",
		X"50",X"E8",X"C8",X"D0",X"E2",X"8D",X"2B",X"18",X"AD",X"28",X"18",X"29",X"03",X"D0",X"06",X"A9",
		X"04",X"8D",X"41",X"03",X"60",X"CE",X"41",X"03",X"D0",X"FA",X"AE",X"42",X"03",X"BC",X"3D",X"03",
		X"4A",X"90",X"0A",X"88",X"88",X"C0",X"16",X"B0",X"0C",X"A0",X"4A",X"D0",X"08",X"C8",X"C8",X"C0",
		X"4C",X"90",X"02",X"A0",X"16",X"98",X"9D",X"3D",X"03",X"D0",X"D4",X"20",X"2E",X"6D",X"A2",X"1A",
		X"20",X"98",X"6C",X"20",X"6A",X"7A",X"A0",X"00",X"8C",X"40",X"03",X"A9",X"E0",X"A2",X"1E",X"8E",
		X"71",X"03",X"20",X"8E",X"7A",X"AE",X"40",X"03",X"BD",X"00",X"03",X"85",X"0A",X"1D",X"01",X"03",
		X"F0",X"7B",X"BD",X"01",X"03",X"85",X"0B",X"A9",X"0A",X"20",X"9E",X"7B",X"A2",X"1C",X"20",X"98",
		X"6C",X"AE",X"40",X"03",X"BD",X"1E",X"03",X"20",X"6A",X"55",X"AE",X"40",X"03",X"BD",X"1F",X"03",
		X"20",X"6A",X"55",X"AE",X"40",X"03",X"BD",X"20",X"03",X"20",X"6A",X"55",X"A0",X"00",X"AE",X"40",
		X"03",X"BD",X"01",X"03",X"F0",X"24",X"AA",X"AD",X"F0",X"33",X"91",X"02",X"C8",X"AD",X"F1",X"33",
		X"91",X"02",X"E0",X"0A",X"90",X"02",X"A2",X"0A",X"C8",X"AD",X"90",X"35",X"91",X"02",X"C8",X"AD",
		X"91",X"35",X"91",X"02",X"CA",X"D0",X"F1",X"20",X"76",X"7A",X"AE",X"40",X"03",X"E0",X"1B",X"B0",
		X"1C",X"E8",X"E8",X"E8",X"8E",X"40",X"03",X"20",X"6A",X"7A",X"AD",X"71",X"03",X"38",X"E9",X"0A",
		X"8D",X"71",X"03",X"AA",X"A9",X"E0",X"A0",X"00",X"4C",X"B2",X"54",X"45",X"52",X"AD",X"00",X"0A",
		X"4A",X"4A",X"4A",X"4A",X"29",X"03",X"F0",X"1C",X"AA",X"BD",X"86",X"38",X"18",X"F8",X"69",X"01",
		X"D8",X"85",X"13",X"A2",X"2A",X"20",X"98",X"6C",X"A9",X"13",X"A0",X"01",X"20",X"A0",X"7B",X"A2",
		X"2C",X"20",X"98",X"6C",X"20",X"74",X"55",X"4C",X"00",X"50",X"A8",X"BE",X"F1",X"33",X"B9",X"F0",
		X"33",X"4C",X"6E",X"7A",X"20",X"1D",X"7A",X"A9",X"00",X"85",X"28",X"24",X"CE",X"10",X"0F",X"AD",
		X"EC",X"02",X"30",X"0A",X"C9",X"04",X"90",X"06",X"AD",X"70",X"03",X"8D",X"00",X"20",X"60",X"48",
		X"8A",X"BA",X"30",X"0B",X"48",X"E6",X"3A",X"A5",X"3A",X"29",X"0F",X"D0",X"04",X"E6",X"39",X"30",
		X"FE",X"98",X"48",X"D8",X"8D",X"00",X"14",X"AD",X"00",X"0C",X"85",X"EB",X"20",X"C3",X"56",X"A5",
		X"E0",X"2A",X"A5",X"E1",X"2A",X"2A",X"48",X"A5",X"E2",X"2A",X"68",X"2A",X"8D",X"00",X"10",X"20",
		X"B9",X"79",X"2C",X"45",X"03",X"30",X"1D",X"A5",X"EF",X"D0",X"19",X"A5",X"D4",X"F0",X"04",X"A9",
		X"20",X"D0",X"0E",X"A5",X"C8",X"F0",X"04",X"A9",X"04",X"D0",X"06",X"24",X"DE",X"10",X"05",X"A9",
		X"40",X"20",X"85",X"79",X"A5",X"0F",X"F0",X"0A",X"C6",X"0F",X"D0",X"04",X"A9",X"00",X"F0",X"02",
		X"A9",X"01",X"A8",X"A5",X"BD",X"F0",X"08",X"C6",X"BD",X"F0",X"04",X"98",X"09",X"04",X"A8",X"98",
		X"05",X"15",X"24",X"CE",X"10",X"05",X"09",X"A0",X"4C",X"94",X"56",X"24",X"CD",X"30",X"7E",X"A9",
		X"00",X"A6",X"EA",X"F0",X"0D",X"09",X"20",X"A6",X"EF",X"D0",X"07",X"48",X"A9",X"20",X"20",X"85",
		X"79",X"68",X"48",X"A5",X"EB",X"29",X"03",X"F0",X"04",X"A5",X"0E",X"F0",X"64",X"A5",X"C6",X"4A",
		X"4A",X"68",X"90",X"02",X"09",X"40",X"8D",X"2B",X"18",X"8D",X"40",X"18",X"AD",X"28",X"18",X"29",
		X"20",X"F0",X"54",X"A9",X"FF",X"8D",X"EC",X"02",X"85",X"CE",X"A5",X"0E",X"38",X"ED",X"70",X"03",
		X"85",X"0E",X"A9",X"00",X"8D",X"2F",X"18",X"85",X"EC",X"8D",X"4B",X"03",X"8D",X"40",X"18",X"85",
		X"B8",X"85",X"B9",X"85",X"BB",X"85",X"BA",X"85",X"C4",X"85",X"26",X"85",X"CD",X"85",X"D2",X"85",
		X"D4",X"85",X"DE",X"85",X"2A",X"85",X"2E",X"85",X"32",X"A9",X"07",X"8D",X"2F",X"18",X"20",X"BE",
		X"69",X"18",X"AD",X"00",X"0A",X"29",X"03",X"69",X"02",X"85",X"CC",X"10",X"0A",X"09",X"60",X"D0",
		X"03",X"68",X"09",X"40",X"8D",X"40",X"18",X"C6",X"ED",X"D0",X"22",X"8D",X"00",X"16",X"A5",X"28",
		X"D0",X"14",X"AD",X"01",X"20",X"49",X"04",X"8D",X"01",X"20",X"29",X"04",X"D0",X"04",X"A9",X"28",
		X"D0",X"02",X"A9",X"20",X"85",X"28",X"8D",X"00",X"12",X"A9",X"06",X"85",X"ED",X"68",X"A8",X"68",
		X"AA",X"68",X"40",X"A2",X"02",X"AD",X"00",X"08",X"E0",X"01",X"F0",X"03",X"B0",X"02",X"4A",X"4A",
		X"4A",X"B5",X"E7",X"29",X"1F",X"B0",X"37",X"F0",X"10",X"C9",X"1B",X"B0",X"0A",X"A8",X"A5",X"3A",
		X"29",X"07",X"C9",X"07",X"98",X"90",X"02",X"E9",X"01",X"95",X"E7",X"AD",X"00",X"08",X"29",X"08",
		X"D0",X"04",X"A9",X"F0",X"85",X"EA",X"A5",X"EA",X"F0",X"08",X"C6",X"EA",X"A9",X"00",X"95",X"E7",
		X"95",X"E4",X"18",X"B5",X"E4",X"F0",X"23",X"D6",X"E4",X"D0",X"1F",X"38",X"B0",X"1C",X"C9",X"1B",
		X"B0",X"09",X"B5",X"E7",X"69",X"20",X"90",X"D1",X"F0",X"01",X"18",X"A9",X"1F",X"B0",X"CA",X"95",
		X"E7",X"B5",X"E4",X"F0",X"01",X"38",X"A9",X"78",X"95",X"E4",X"90",X"2A",X"A9",X"00",X"E0",X"01",
		X"90",X"16",X"F0",X"0C",X"A5",X"EB",X"29",X"0C",X"4A",X"4A",X"F0",X"0C",X"69",X"02",X"D0",X"08",
		X"A5",X"EB",X"29",X"10",X"F0",X"02",X"A9",X"01",X"38",X"48",X"65",X"EC",X"85",X"EC",X"68",X"38",
		X"65",X"21",X"85",X"21",X"F6",X"E0",X"CA",X"30",X"03",X"4C",X"C5",X"56",X"A5",X"EB",X"4A",X"4A",
		X"4A",X"4A",X"4A",X"A8",X"A5",X"EC",X"38",X"F9",X"78",X"57",X"30",X"14",X"85",X"EC",X"E6",X"21",
		X"C0",X"03",X"D0",X"0C",X"E6",X"21",X"D0",X"08",X"7F",X"02",X"04",X"04",X"05",X"7F",X"7F",X"7F",
		X"A5",X"EB",X"29",X"03",X"A8",X"F0",X"12",X"4A",X"69",X"00",X"49",X"FF",X"38",X"65",X"21",X"90",
		X"0A",X"C0",X"02",X"B0",X"02",X"E6",X"0E",X"E6",X"0E",X"85",X"21",X"A5",X"3A",X"4A",X"B0",X"27",
		X"A0",X"00",X"A2",X"02",X"B5",X"E0",X"F0",X"09",X"C9",X"10",X"90",X"05",X"69",X"EF",X"C8",X"95",
		X"E0",X"CA",X"10",X"F0",X"98",X"D0",X"10",X"A2",X"02",X"B5",X"E0",X"F0",X"07",X"18",X"69",X"EF",
		X"95",X"E0",X"30",X"03",X"CA",X"10",X"F2",X"60",X"A2",X"00",X"86",X"07",X"86",X"06",X"A5",X"27",
		X"85",X"04",X"A5",X"2A",X"4A",X"66",X"04",X"4A",X"66",X"04",X"4A",X"66",X"04",X"4A",X"66",X"04",
		X"48",X"29",X"01",X"09",X"02",X"85",X"05",X"A5",X"DF",X"4A",X"4A",X"4A",X"4A",X"F0",X"0D",X"85",
		X"08",X"38",X"A5",X"06",X"E5",X"08",X"85",X"06",X"A9",X"FF",X"85",X"07",X"20",X"6A",X"7A",X"20",
		X"AB",X"7A",X"A9",X"30",X"A2",X"00",X"20",X"5A",X"7A",X"68",X"49",X"0F",X"20",X"A7",X"58",X"20",
		X"A7",X"58",X"20",X"A7",X"58",X"A5",X"27",X"85",X"04",X"A5",X"2A",X"C9",X"88",X"B0",X"04",X"C9",
		X"39",X"B0",X"01",X"60",X"4A",X"66",X"04",X"4A",X"66",X"04",X"4A",X"66",X"04",X"4A",X"66",X"04",
		X"85",X"05",X"A5",X"04",X"38",X"E9",X"05",X"85",X"04",X"A5",X"05",X"E9",X"06",X"85",X"05",X"18",
		X"A9",X"5E",X"65",X"06",X"85",X"06",X"90",X"02",X"E6",X"07",X"20",X"6A",X"7A",X"20",X"AB",X"7A",
		X"A9",X"00",X"85",X"35",X"85",X"36",X"85",X"37",X"85",X"38",X"A2",X"04",X"BD",X"4D",X"03",X"F0",
		X"42",X"BD",X"5C",X"03",X"38",X"A8",X"E5",X"35",X"85",X"04",X"84",X"35",X"BD",X"61",X"03",X"A8",
		X"E5",X"36",X"85",X"05",X"84",X"36",X"38",X"BD",X"66",X"03",X"A8",X"E5",X"37",X"85",X"06",X"84",
		X"37",X"BD",X"6B",X"03",X"A8",X"E5",X"38",X"85",X"07",X"84",X"38",X"A9",X"00",X"85",X"01",X"86",
		X"08",X"20",X"AB",X"7A",X"A6",X"08",X"BD",X"4D",X"03",X"0A",X"0A",X"0A",X"29",X"E0",X"20",X"8A",
		X"7A",X"A6",X"08",X"CA",X"10",X"B6",X"60",X"29",X"0E",X"A8",X"B9",X"06",X"30",X"C8",X"BE",X"06",
		X"30",X"C8",X"84",X"08",X"20",X"6E",X"7A",X"A5",X"08",X"60",X"A2",X"04",X"BD",X"4D",X"03",X"D0",
		X"37",X"AD",X"2A",X"18",X"29",X"07",X"D0",X"77",X"A9",X"1F",X"9D",X"4D",X"03",X"AD",X"2A",X"18",
		X"29",X"03",X"69",X"01",X"2C",X"2A",X"18",X"50",X"02",X"49",X"FF",X"9D",X"52",X"03",X"AD",X"2A",
		X"18",X"29",X"07",X"69",X"05",X"9D",X"57",X"03",X"A9",X"00",X"9D",X"5C",X"03",X"9D",X"61",X"03",
		X"9D",X"66",X"03",X"9D",X"6B",X"03",X"F0",X"47",X"DE",X"4D",X"03",X"F0",X"EB",X"DE",X"57",X"03",
		X"A0",X"00",X"18",X"BD",X"57",X"03",X"10",X"01",X"88",X"7D",X"66",X"03",X"9D",X"66",X"03",X"BD",
		X"6B",X"03",X"10",X"0E",X"BD",X"66",X"03",X"C9",X"A2",X"B0",X"07",X"A9",X"00",X"9D",X"4D",X"03",
		X"F0",X"C6",X"98",X"7D",X"6B",X"03",X"9D",X"6B",X"03",X"A0",X"00",X"18",X"BD",X"52",X"03",X"10",
		X"01",X"88",X"7D",X"5C",X"03",X"9D",X"5C",X"03",X"98",X"7D",X"61",X"03",X"9D",X"61",X"03",X"CA",
		X"30",X"03",X"4C",X"BC",X"58",X"60",X"A0",X"00",X"A5",X"2D",X"8D",X"64",X"18",X"A5",X"2E",X"8D",
		X"65",X"18",X"A5",X"31",X"8D",X"66",X"18",X"A5",X"32",X"8D",X"67",X"18",X"A5",X"27",X"18",X"2A",
		X"2A",X"A6",X"2A",X"20",X"17",X"5F",X"49",X"FF",X"69",X"01",X"8D",X"62",X"18",X"8A",X"49",X"FF",
		X"69",X"00",X"8D",X"63",X"18",X"A5",X"A6",X"A6",X"2A",X"20",X"F9",X"5E",X"8D",X"60",X"18",X"8E",
		X"61",X"18",X"2C",X"4B",X"03",X"10",X"05",X"A2",X"00",X"4C",X"EE",X"5A",X"A5",X"14",X"F0",X"06",
		X"20",X"89",X"5B",X"4C",X"6C",X"5A",X"A5",X"2C",X"8D",X"71",X"02",X"A9",X"16",X"24",X"CB",X"30",
		X"0A",X"A2",X"21",X"20",X"B5",X"69",X"B0",X"02",X"A2",X"02",X"8A",X"8D",X"70",X"02",X"A5",X"2F",
		X"8D",X"68",X"18",X"A5",X"30",X"8D",X"69",X"18",X"A5",X"33",X"8D",X"6A",X"18",X"A5",X"34",X"8D",
		X"6B",X"18",X"20",X"1F",X"5B",X"98",X"F0",X"CB",X"AD",X"71",X"02",X"99",X"71",X"02",X"AD",X"00",
		X"02",X"99",X"00",X"02",X"AD",X"01",X"02",X"99",X"01",X"02",X"AD",X"38",X"02",X"99",X"38",X"02",
		X"AD",X"39",X"02",X"99",X"39",X"02",X"24",X"CB",X"10",X"09",X"A5",X"A7",X"29",X"07",X"18",X"69",
		X"24",X"D0",X"1D",X"20",X"B5",X"69",X"B0",X"74",X"AD",X"71",X"02",X"38",X"E5",X"2A",X"18",X"69",
		X"40",X"0A",X"A9",X"04",X"90",X"01",X"0A",X"85",X"08",X"A5",X"A7",X"29",X"03",X"18",X"65",X"08",
		X"99",X"70",X"02",X"C8",X"C8",X"24",X"CB",X"30",X"53",X"A9",X"0D",X"99",X"70",X"02",X"A5",X"BE",
		X"99",X"71",X"02",X"A5",X"2A",X"38",X"E5",X"2C",X"85",X"2B",X"20",X"4B",X"5E",X"8A",X"A2",X"FF",
		X"49",X"FF",X"30",X"01",X"E8",X"18",X"69",X"01",X"90",X"01",X"E8",X"0A",X"48",X"8A",X"2A",X"AA",
		X"68",X"18",X"6D",X"00",X"02",X"99",X"00",X"02",X"8A",X"6D",X"01",X"02",X"99",X"01",X"02",X"A5",
		X"2B",X"20",X"4E",X"5E",X"8A",X"0A",X"A2",X"00",X"90",X"02",X"A2",X"FF",X"18",X"6D",X"38",X"02",
		X"99",X"38",X"02",X"8A",X"6D",X"39",X"02",X"99",X"39",X"02",X"C8",X"C8",X"A2",X"02",X"B5",X"24",
		X"F0",X"40",X"B5",X"2A",X"99",X"71",X"02",X"A9",X"03",X"99",X"70",X"02",X"B5",X"24",X"10",X"1B",
		X"18",X"69",X"0F",X"30",X"06",X"A9",X"00",X"95",X"24",X"F0",X"27",X"95",X"24",X"49",X"FF",X"18",
		X"79",X"01",X"02",X"99",X"71",X"02",X"A9",X"0E",X"99",X"70",X"02",X"B5",X"A8",X"8D",X"68",X"18",
		X"B5",X"A9",X"8D",X"69",X"18",X"B5",X"AC",X"8D",X"6A",X"18",X"B5",X"AD",X"8D",X"6B",X"18",X"20",
		X"1F",X"5B",X"CA",X"CA",X"10",X"B8",X"A5",X"DE",X"F0",X"32",X"A9",X"20",X"99",X"70",X"02",X"A5",
		X"D9",X"99",X"71",X"02",X"A5",X"D5",X"8D",X"68",X"18",X"A5",X"D6",X"8D",X"69",X"18",X"A5",X"D7",
		X"8D",X"6A",X"18",X"A5",X"D8",X"8D",X"6B",X"18",X"20",X"1F",X"5B",X"B9",X"6E",X"02",X"C9",X"20",
		X"D0",X"06",X"A9",X"81",X"85",X"DE",X"D0",X"04",X"A9",X"01",X"85",X"DE",X"A2",X"00",X"BD",X"CC",
		X"3F",X"30",X"28",X"99",X"70",X"02",X"BD",X"CD",X"3F",X"99",X"71",X"02",X"BD",X"81",X"76",X"8D",
		X"68",X"18",X"BD",X"82",X"76",X"8D",X"69",X"18",X"BD",X"AB",X"76",X"8D",X"6A",X"18",X"BD",X"AC",
		X"76",X"8D",X"6B",X"18",X"20",X"1F",X"5B",X"E8",X"E8",X"D0",X"D3",X"99",X"70",X"02",X"60",X"20",
		X"80",X"5B",X"0A",X"85",X"1B",X"AD",X"18",X"18",X"8D",X"72",X"18",X"30",X"52",X"2A",X"30",X"4F",
		X"85",X"1C",X"4A",X"4A",X"F0",X"49",X"A5",X"1C",X"C9",X"7B",X"B0",X"43",X"20",X"80",X"5B",X"0A",
		X"85",X"1F",X"AD",X"18",X"18",X"2A",X"85",X"20",X"A5",X"1F",X"24",X"20",X"10",X"05",X"18",X"49",
		X"FF",X"69",X"01",X"85",X"1D",X"A5",X"20",X"10",X"04",X"49",X"FF",X"69",X"00",X"85",X"1E",X"A5",
		X"1D",X"C5",X"1B",X"A5",X"1E",X"E5",X"1C",X"B0",X"16",X"A5",X"1B",X"99",X"00",X"02",X"A5",X"1C",
		X"99",X"01",X"02",X"A5",X"1F",X"99",X"38",X"02",X"A5",X"20",X"99",X"39",X"02",X"C8",X"C8",X"60",
		X"2C",X"00",X"18",X"30",X"FB",X"AD",X"10",X"18",X"60",X"A2",X"0A",X"BD",X"D9",X"02",X"18",X"10",
		X"03",X"4C",X"3D",X"5C",X"BD",X"A8",X"02",X"7D",X"AE",X"3F",X"9D",X"A8",X"02",X"8D",X"68",X"18",
		X"BD",X"A9",X"02",X"7D",X"AF",X"3F",X"9D",X"A9",X"02",X"8D",X"69",X"18",X"18",X"BD",X"B8",X"02",
		X"7D",X"BA",X"3F",X"9D",X"B8",X"02",X"8D",X"6A",X"18",X"BD",X"B9",X"02",X"7D",X"BB",X"3F",X"9D",
		X"B9",X"02",X"BD",X"C9",X"02",X"85",X"08",X"30",X"02",X"A9",X"00",X"F0",X"02",X"A9",X"FF",X"06",
		X"08",X"2A",X"06",X"08",X"2A",X"85",X"09",X"BD",X"D8",X"02",X"18",X"65",X"08",X"9D",X"D8",X"02",
		X"A5",X"09",X"7D",X"D9",X"02",X"9D",X"D9",X"02",X"BD",X"C9",X"02",X"10",X"04",X"C9",X"85",X"90",
		X"05",X"69",X"FC",X"9D",X"C9",X"02",X"8A",X"4A",X"4A",X"08",X"8A",X"0A",X"0A",X"69",X"03",X"28",
		X"90",X"0A",X"85",X"08",X"BD",X"C8",X"02",X"E5",X"08",X"4C",X"0F",X"5C",X"7D",X"C8",X"02",X"9D",
		X"C8",X"02",X"99",X"71",X"02",X"8A",X"4A",X"18",X"69",X"10",X"24",X"CB",X"10",X"04",X"69",X"08",
		X"D0",X"0F",X"C9",X"13",X"D0",X"0B",X"85",X"08",X"20",X"B5",X"69",X"90",X"02",X"E6",X"08",X"A5",
		X"08",X"99",X"70",X"02",X"BD",X"B9",X"02",X"8D",X"6B",X"18",X"20",X"1F",X"5B",X"CA",X"CA",X"30",
		X"03",X"4C",X"8B",X"5B",X"A2",X"0A",X"BD",X"D9",X"02",X"10",X"0F",X"CA",X"CA",X"10",X"F7",X"A9",
		X"00",X"85",X"14",X"98",X"48",X"20",X"BE",X"69",X"68",X"A8",X"60",X"5E",X"0A",X"A8",X"B9",X"72",
		X"74",X"85",X"3B",X"B9",X"73",X"74",X"85",X"3C",X"A0",X"00",X"B1",X"3B",X"C9",X"FF",X"D0",X"01",
		X"60",X"AA",X"29",X"F8",X"85",X"08",X"8A",X"29",X"07",X"0A",X"AA",X"BD",X"85",X"5C",X"48",X"BD",
		X"84",X"5C",X"48",X"60",X"91",X"5C",X"9E",X"5C",X"E0",X"5C",X"D3",X"5C",X"E4",X"5C",X"EC",X"5C",
		X"0D",X"5D",X"A9",X"00",X"20",X"11",X"5D",X"A9",X"20",X"20",X"8A",X"7A",X"4C",X"41",X"5D",X"A6",
		X"10",X"BD",X"70",X"02",X"C9",X"17",X"F0",X"10",X"C9",X"1E",X"F0",X"0C",X"C9",X"1F",X"F0",X"08",
		X"C9",X"20",X"D0",X"0A",X"A5",X"D4",X"F0",X"06",X"AD",X"EA",X"02",X"4C",X"CB",X"5C",X"A5",X"08",
		X"38",X"E5",X"25",X"90",X"04",X"C9",X"30",X"B0",X"02",X"A9",X"30",X"A8",X"A9",X"04",X"20",X"63",
		X"7A",X"4C",X"41",X"5D",X"A9",X"00",X"85",X"35",X"85",X"36",X"85",X"37",X"85",X"38",X"20",X"6A",
		X"7A",X"A9",X"00",X"F0",X"02",X"A9",X"20",X"20",X"11",X"5D",X"4C",X"41",X"5D",X"A6",X"10",X"BD",
		X"71",X"02",X"AA",X"29",X"3F",X"0A",X"A8",X"8A",X"29",X"C0",X"0A",X"2A",X"2A",X"69",X"01",X"20",
		X"83",X"7A",X"A2",X"7A",X"A9",X"34",X"20",X"5A",X"7A",X"A9",X"01",X"20",X"81",X"7A",X"4C",X"41",
		X"5D",X"85",X"01",X"A5",X"08",X"4A",X"AA",X"B5",X"3D",X"A8",X"38",X"E5",X"35",X"85",X"04",X"84",
		X"35",X"B5",X"3E",X"A8",X"E5",X"36",X"85",X"05",X"84",X"36",X"38",X"B5",X"3F",X"A8",X"E5",X"37",
		X"85",X"06",X"84",X"37",X"B5",X"40",X"A8",X"E5",X"38",X"85",X"07",X"84",X"38",X"20",X"AB",X"7A",
		X"60",X"E6",X"3B",X"D0",X"02",X"E6",X"3C",X"4C",X"68",X"5C",X"86",X"13",X"A5",X"2A",X"38",X"FD",
		X"71",X"02",X"49",X"80",X"85",X"2B",X"20",X"4E",X"5E",X"8D",X"62",X"18",X"8E",X"63",X"18",X"A5",
		X"2B",X"20",X"4B",X"5E",X"18",X"49",X"FF",X"69",X"01",X"8D",X"60",X"18",X"8A",X"49",X"FF",X"69",
		X"00",X"8D",X"61",X"18",X"A6",X"13",X"BD",X"70",X"02",X"0A",X"A8",X"B9",X"8E",X"38",X"85",X"3B",
		X"B9",X"8F",X"38",X"85",X"3C",X"BD",X"00",X"02",X"8D",X"64",X"18",X"BD",X"01",X"02",X"8D",X"65",
		X"18",X"29",X"F0",X"85",X"25",X"BD",X"38",X"02",X"8D",X"66",X"18",X"BD",X"39",X"02",X"8D",X"67",
		X"18",X"A2",X"00",X"8E",X"6D",X"18",X"8E",X"6E",X"18",X"86",X"18",X"E6",X"18",X"A4",X"18",X"B1",
		X"3B",X"8D",X"68",X"18",X"C8",X"B1",X"3B",X"8D",X"69",X"18",X"C8",X"B1",X"3B",X"8D",X"6A",X"18",
		X"C8",X"B1",X"3B",X"8D",X"71",X"18",X"C8",X"20",X"80",X"5B",X"18",X"49",X"FF",X"69",X"01",X"95",
		X"3D",X"AD",X"18",X"18",X"49",X"FF",X"69",X"00",X"95",X"3E",X"B1",X"3B",X"85",X"22",X"C8",X"B1",
		X"3B",X"C8",X"84",X"18",X"85",X"23",X"86",X"16",X"20",X"05",X"5E",X"20",X"80",X"5B",X"A6",X"16",
		X"95",X"3F",X"AD",X"18",X"18",X"95",X"40",X"98",X"A0",X"00",X"D1",X"3B",X"B0",X"06",X"E8",X"E8",
		X"E8",X"E8",X"D0",X"A9",X"60",X"A6",X"13",X"BD",X"70",X"02",X"29",X"10",X"F0",X"15",X"BD",X"70",
		X"02",X"29",X"07",X"0A",X"AA",X"BD",X"D8",X"02",X"65",X"22",X"85",X"22",X"BD",X"D9",X"02",X"65",
		X"23",X"85",X"23",X"A5",X"DF",X"F0",X"0F",X"38",X"A5",X"22",X"E5",X"DF",X"8D",X"6F",X"18",X"A5",
		X"23",X"E9",X"00",X"4C",X"3D",X"5E",X"A5",X"22",X"8D",X"6F",X"18",X"A5",X"23",X"8D",X"70",X"18",
		X"8D",X"74",X"18",X"60",X"A5",X"DF",X"F0",X"02",X"46",X"DF",X"60",X"18",X"69",X"40",X"10",X"13",
		X"29",X"7F",X"20",X"63",X"5E",X"49",X"FF",X"18",X"69",X"01",X"48",X"8A",X"49",X"FF",X"69",X"00",
		X"AA",X"68",X"60",X"C9",X"41",X"90",X"04",X"49",X"7F",X"69",X"00",X"0A",X"AA",X"BD",X"77",X"5E",
		X"48",X"BD",X"78",X"5E",X"AA",X"68",X"60",X"00",X"00",X"24",X"03",X"47",X"06",X"6A",X"09",X"8B",
		X"0C",X"AB",X"0F",X"C8",X"12",X"E2",X"15",X"F8",X"18",X"0B",X"1C",X"19",X"1F",X"23",X"22",X"28",
		X"25",X"26",X"28",X"1F",X"2B",X"11",X"2E",X"FB",X"30",X"DE",X"33",X"BE",X"36",X"8C",X"39",X"56",
		X"3C",X"17",X"3F",X"CE",X"41",X"7A",X"44",X"1C",X"47",X"B4",X"49",X"3F",X"4C",X"BF",X"4E",X"33",
		X"51",X"9B",X"53",X"F5",X"55",X"42",X"58",X"82",X"5A",X"B4",X"5C",X"D7",X"5E",X"EC",X"60",X"F2",
		X"62",X"EB",X"64",X"CF",X"66",X"A6",X"68",X"6D",X"6A",X"24",X"6C",X"C4",X"6D",X"5F",X"6F",X"E2",
		X"70",X"55",X"72",X"B5",X"73",X"04",X"75",X"41",X"76",X"6C",X"77",X"84",X"78",X"8A",X"79",X"7D",
		X"7A",X"5D",X"7B",X"2A",X"7C",X"E3",X"7C",X"8A",X"7D",X"1D",X"7E",X"9D",X"7E",X"09",X"7F",X"62",
		X"7F",X"A7",X"7F",X"D8",X"7F",X"F6",X"7F",X"FF",X"7F",X"29",X"01",X"85",X"A6",X"D0",X"04",X"8A",
		X"4C",X"4B",X"5E",X"8A",X"85",X"0C",X"20",X"4B",X"5E",X"85",X"08",X"86",X"09",X"E6",X"0C",X"A5",
		X"0C",X"20",X"4B",X"5E",X"4C",X"32",X"5F",X"29",X"01",X"85",X"A6",X"D0",X"04",X"8A",X"4C",X"4E",
		X"5E",X"8A",X"85",X"0C",X"20",X"4E",X"5E",X"85",X"08",X"86",X"09",X"E6",X"0C",X"A5",X"0C",X"20",
		X"4E",X"5E",X"38",X"E5",X"08",X"85",X"0A",X"8A",X"E5",X"09",X"C9",X"80",X"6A",X"66",X"0A",X"85",
		X"0B",X"A5",X"08",X"18",X"65",X"0A",X"48",X"A5",X"09",X"65",X"0B",X"AA",X"68",X"60",X"A5",X"24",
		X"30",X"02",X"D0",X"03",X"4C",X"43",X"60",X"A2",X"00",X"A0",X"02",X"B5",X"A8",X"8D",X"60",X"18",
		X"B5",X"A9",X"8D",X"61",X"18",X"B5",X"AC",X"8D",X"62",X"18",X"B5",X"AD",X"8D",X"63",X"18",X"B9",
		X"12",X"00",X"D0",X"2A",X"B9",X"2D",X"00",X"8D",X"64",X"18",X"B9",X"2E",X"00",X"8D",X"65",X"18",
		X"B9",X"31",X"00",X"8D",X"66",X"18",X"B9",X"32",X"00",X"8D",X"7D",X"18",X"C1",X"00",X"B1",X"00",
		X"AD",X"10",X"18",X"85",X"0C",X"AD",X"18",X"18",X"30",X"3F",X"4A",X"66",X"0C",X"4A",X"D0",X"39",
		X"66",X"0C",X"24",X"CB",X"10",X"0C",X"AD",X"E4",X"02",X"C9",X"00",X"AD",X"E5",X"02",X"E9",X"02",
		X"B0",X"27",X"A5",X"2A",X"38",X"E5",X"2C",X"0A",X"10",X"05",X"49",X"FF",X"18",X"69",X"01",X"4A",
		X"4A",X"24",X"CB",X"30",X"03",X"4A",X"10",X"03",X"18",X"69",X"18",X"85",X"08",X"4A",X"18",X"65",
		X"08",X"69",X"38",X"85",X"08",X"C5",X"0C",X"B0",X"03",X"4C",X"43",X"60",X"A9",X"20",X"99",X"12",
		X"00",X"A9",X"00",X"85",X"D2",X"98",X"D0",X"0E",X"A9",X"02",X"85",X"C7",X"A9",X"FF",X"85",X"DF",
		X"C6",X"CC",X"D0",X"02",X"E6",X"CD",X"B5",X"B8",X"85",X"08",X"B5",X"B9",X"85",X"09",X"8A",X"D0",
		X"0D",X"A9",X"02",X"24",X"CB",X"30",X"09",X"20",X"B5",X"69",X"A9",X"03",X"B0",X"02",X"A9",X"01",
		X"18",X"F8",X"75",X"B8",X"95",X"B8",X"B5",X"B9",X"69",X"00",X"D8",X"95",X"B9",X"8A",X"D0",X"03",
		X"20",X"5F",X"61",X"A9",X"80",X"95",X"24",X"A9",X"FF",X"99",X"0F",X"00",X"A9",X"02",X"19",X"15",
		X"00",X"99",X"15",X"00",X"B5",X"15",X"29",X"FD",X"95",X"15",X"20",X"99",X"61",X"A9",X"70",X"95",
		X"0F",X"38",X"60",X"18",X"60",X"A2",X"02",X"8A",X"49",X"02",X"A8",X"B5",X"24",X"30",X"6B",X"F0",
		X"69",X"A5",X"C7",X"D0",X"04",X"A5",X"CD",X"D0",X"61",X"20",X"5B",X"5F",X"B0",X"5C",X"4C",X"C2",
		X"60",X"A0",X"00",X"B9",X"CC",X"3F",X"30",X"52",X"B9",X"81",X"76",X"8D",X"64",X"18",X"B9",X"82",
		X"76",X"8D",X"65",X"18",X"B9",X"AB",X"76",X"8D",X"66",X"18",X"B9",X"AC",X"76",X"8D",X"7D",X"18",
		X"C1",X"00",X"AD",X"10",X"18",X"85",X"0C",X"AD",X"18",X"18",X"C9",X"80",X"6A",X"66",X"0C",X"C9",
		X"80",X"6A",X"66",X"0C",X"C9",X"00",X"D0",X"1E",X"86",X"A6",X"BE",X"CC",X"3F",X"BD",X"39",X"61",
		X"A6",X"A6",X"C5",X"0C",X"90",X"10",X"A9",X"A0",X"95",X"24",X"A9",X"70",X"85",X"0F",X"A5",X"15",
		X"29",X"FD",X"85",X"15",X"B0",X"04",X"C8",X"C8",X"D0",X"A9",X"CA",X"CA",X"D0",X"03",X"4C",X"47",
		X"60",X"60",X"A5",X"DE",X"F0",X"33",X"A5",X"D4",X"D0",X"2F",X"A5",X"D5",X"8D",X"64",X"18",X"A5",
		X"D6",X"8D",X"65",X"18",X"A5",X"D7",X"8D",X"66",X"18",X"A5",X"D8",X"8D",X"67",X"18",X"8D",X"7D",
		X"18",X"C1",X"00",X"AD",X"10",X"18",X"85",X"0C",X"AD",X"18",X"18",X"C9",X"80",X"6A",X"66",X"0C",
		X"C9",X"80",X"6A",X"66",X"0C",X"C9",X"00",X"F0",X"03",X"4C",X"61",X"60",X"A9",X"90",X"C5",X"0C",
		X"90",X"F7",X"A9",X"40",X"85",X"D4",X"A9",X"20",X"20",X"85",X"79",X"A9",X"A0",X"95",X"24",X"95",
		X"0F",X"A9",X"02",X"19",X"15",X"00",X"99",X"15",X"00",X"8A",X"D0",X"9E",X"A5",X"B8",X"85",X"08",
		X"A5",X"B9",X"85",X"09",X"A9",X"05",X"18",X"F8",X"65",X"B8",X"85",X"B8",X"A5",X"B9",X"69",X"00",
		X"D8",X"85",X"B9",X"20",X"5F",X"61",X"4C",X"BA",X"60",X"38",X"58",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"56",X"00",X"00",X"00",X"24",X"09",X"10",X"11",X"A5",X"08",X"18",
		X"49",X"FF",X"69",X"01",X"85",X"08",X"A5",X"09",X"49",X"FF",X"69",X"00",X"85",X"09",X"60",X"AD",
		X"00",X"0A",X"4A",X"4A",X"4A",X"4A",X"29",X"03",X"AA",X"BD",X"86",X"38",X"F0",X"17",X"A6",X"B9",
		X"D0",X"16",X"C5",X"08",X"90",X"0F",X"C5",X"B8",X"B0",X"0B",X"E6",X"CC",X"A9",X"00",X"85",X"CD",
		X"A9",X"08",X"20",X"85",X"79",X"A2",X"00",X"60",X"A5",X"09",X"D0",X"F9",X"85",X"CD",X"E6",X"CC",
		X"A9",X"FF",X"8D",X"45",X"03",X"A9",X"80",X"D0",X"E9",X"8A",X"D0",X"33",X"A2",X"05",X"A0",X"0A",
		X"BD",X"C6",X"3F",X"99",X"C9",X"02",X"A5",X"2F",X"99",X"A8",X"02",X"A5",X"30",X"99",X"A9",X"02",
		X"A5",X"33",X"99",X"B8",X"02",X"A5",X"34",X"99",X"B9",X"02",X"AD",X"2A",X"18",X"99",X"C8",X"02",
		X"A9",X"00",X"99",X"D8",X"02",X"99",X"D9",X"02",X"88",X"88",X"CA",X"10",X"D3",X"A2",X"00",X"60",
		X"24",X"CE",X"30",X"24",X"2C",X"4B",X"03",X"30",X"25",X"A5",X"C7",X"D0",X"21",X"A2",X"00",X"24",
		X"C6",X"70",X"06",X"20",X"51",X"63",X"4C",X"EC",X"61",X"20",X"6F",X"63",X"24",X"30",X"10",X"05",
		X"50",X"0C",X"4C",X"8D",X"63",X"4C",X"9B",X"63",X"A2",X"00",X"B5",X"12",X"F0",X"01",X"60",X"20",
		X"A9",X"63",X"8E",X"2B",X"18",X"AD",X"28",X"18",X"8D",X"EB",X"02",X"49",X"0F",X"29",X"0F",X"C9",
		X"05",X"90",X"7F",X"0A",X"A8",X"B9",X"15",X"62",X"48",X"B9",X"14",X"62",X"48",X"60",X"5D",X"62",
		X"33",X"62",X"51",X"62",X"91",X"62",X"3C",X"62",X"68",X"62",X"4B",X"62",X"91",X"62",X"45",X"62",
		X"57",X"62",X"91",X"62",X"20",X"9B",X"63",X"20",X"9B",X"63",X"4C",X"8A",X"62",X"20",X"8D",X"63",
		X"20",X"8D",X"63",X"4C",X"8A",X"62",X"20",X"8D",X"63",X"4C",X"61",X"62",X"20",X"8D",X"63",X"4C",
		X"6C",X"62",X"20",X"9B",X"63",X"4C",X"61",X"62",X"20",X"9B",X"63",X"4C",X"6C",X"62",X"20",X"51",
		X"63",X"20",X"51",X"63",X"F6",X"A5",X"4C",X"71",X"62",X"20",X"6F",X"63",X"20",X"6F",X"63",X"D6",
		X"A5",X"20",X"D6",X"68",X"90",X"14",X"20",X"BA",X"63",X"A5",X"C8",X"D0",X"11",X"A9",X"02",X"20",
		X"85",X"79",X"A9",X"3F",X"85",X"DF",X"E6",X"C8",X"D0",X"04",X"A9",X"00",X"85",X"C8",X"A9",X"10",
		X"D0",X"02",X"A9",X"00",X"85",X"08",X"BD",X"15",X"00",X"29",X"EF",X"05",X"08",X"95",X"15",X"B5",
		X"24",X"D0",X"6C",X"AD",X"EB",X"02",X"29",X"10",X"F0",X"65",X"A9",X"7F",X"95",X"24",X"B5",X"15",
		X"09",X"08",X"95",X"15",X"A9",X"05",X"85",X"BD",X"B5",X"27",X"18",X"2A",X"2A",X"48",X"B5",X"2A",
		X"86",X"13",X"AA",X"68",X"20",X"F9",X"5E",X"85",X"08",X"8A",X"08",X"A6",X"13",X"95",X"B0",X"28",
		X"30",X"04",X"A9",X"00",X"F0",X"02",X"A9",X"FF",X"06",X"08",X"36",X"B0",X"2A",X"95",X"B1",X"B5",
		X"2A",X"AA",X"A5",X"A6",X"20",X"17",X"5F",X"85",X"08",X"8A",X"08",X"A6",X"13",X"95",X"B4",X"28",
		X"30",X"04",X"A9",X"00",X"F0",X"02",X"A9",X"FF",X"06",X"08",X"36",X"B4",X"2A",X"95",X"B5",X"B5",
		X"2D",X"95",X"A8",X"B5",X"2E",X"95",X"A9",X"B5",X"31",X"95",X"AC",X"B5",X"32",X"95",X"AD",X"60",
		X"B5",X"2A",X"86",X"08",X"20",X"4E",X"5E",X"8A",X"C9",X"80",X"6A",X"85",X"1D",X"C9",X"80",X"6A",
		X"18",X"65",X"1D",X"85",X"1D",X"10",X"04",X"A9",X"FF",X"30",X"02",X"A9",X"00",X"85",X"1E",X"A6",
		X"08",X"B5",X"2A",X"20",X"4B",X"5E",X"8A",X"C9",X"80",X"6A",X"85",X"19",X"C9",X"80",X"6A",X"18",
		X"65",X"19",X"85",X"19",X"10",X"04",X"A9",X"FF",X"30",X"02",X"A9",X"00",X"85",X"1A",X"A6",X"08",
		X"60",X"20",X"10",X"63",X"B5",X"2D",X"18",X"65",X"19",X"95",X"2D",X"B5",X"2E",X"65",X"1A",X"95",
		X"2E",X"B5",X"31",X"18",X"65",X"1D",X"95",X"31",X"B5",X"32",X"65",X"1E",X"95",X"32",X"60",X"20",
		X"10",X"63",X"B5",X"2D",X"38",X"E5",X"19",X"95",X"2D",X"B5",X"2E",X"E5",X"1A",X"95",X"2E",X"38",
		X"B5",X"31",X"E5",X"1D",X"95",X"31",X"B5",X"32",X"E5",X"1E",X"95",X"32",X"60",X"A9",X"80",X"18",
		X"75",X"27",X"95",X"27",X"A9",X"00",X"75",X"2A",X"95",X"2A",X"60",X"B5",X"27",X"38",X"E9",X"80",
		X"95",X"27",X"B5",X"2A",X"E9",X"00",X"95",X"2A",X"60",X"B5",X"2D",X"85",X"C0",X"B5",X"2E",X"85",
		X"C1",X"B5",X"31",X"85",X"C2",X"B5",X"32",X"85",X"C3",X"60",X"A5",X"C0",X"95",X"2D",X"A5",X"C1",
		X"95",X"2E",X"A5",X"C2",X"95",X"31",X"A5",X"C3",X"95",X"32",X"60",X"48",X"24",X"CE",X"30",X"1D",
		X"A9",X"30",X"85",X"C4",X"D0",X"3A",X"A5",X"B9",X"F0",X"06",X"A9",X"7F",X"85",X"CF",X"D0",X"1D",
		X"A5",X"B8",X"38",X"E5",X"BA",X"85",X"CF",X"B0",X"04",X"49",X"FF",X"69",X"01",X"C9",X"05",X"B0",
		X"0C",X"85",X"C4",X"A9",X"05",X"E5",X"C4",X"0A",X"0A",X"0A",X"0A",X"D0",X"02",X"A9",X"04",X"85",
		X"C4",X"24",X"CF",X"30",X"0B",X"A9",X"0A",X"38",X"E5",X"CF",X"B0",X"06",X"A9",X"01",X"D0",X"02",
		X"A9",X"0A",X"0A",X"85",X"CF",X"68",X"60",X"D5",X"A5",X"14",X"F0",X"01",X"60",X"24",X"CB",X"10",
		X"03",X"4C",X"24",X"66",X"A2",X"02",X"20",X"A9",X"63",X"18",X"A5",X"BE",X"69",X"0B",X"85",X"BE",
		X"A5",X"C5",X"4A",X"90",X"27",X"4A",X"08",X"20",X"6F",X"63",X"28",X"90",X"06",X"20",X"8D",X"63",
		X"4C",X"46",X"64",X"20",X"9B",X"63",X"C6",X"A7",X"A5",X"C4",X"F0",X"01",X"60",X"A5",X"C5",X"29",
		X"FC",X"85",X"C5",X"A5",X"2C",X"85",X"BC",X"A9",X"34",X"85",X"C4",X"60",X"A5",X"C4",X"D0",X"03",
		X"4C",X"34",X"65",X"A5",X"2C",X"38",X"E5",X"BC",X"A8",X"10",X"05",X"49",X"FF",X"18",X"69",X"01",
		X"C5",X"CF",X"90",X"3E",X"98",X"10",X"1E",X"20",X"8D",X"63",X"20",X"95",X"65",X"20",X"8D",X"63",
		X"20",X"95",X"65",X"20",X"B5",X"69",X"B0",X"01",X"60",X"20",X"8D",X"63",X"20",X"95",X"65",X"20",
		X"8D",X"63",X"4C",X"95",X"65",X"20",X"9B",X"63",X"20",X"95",X"65",X"20",X"9B",X"63",X"20",X"95",
		X"65",X"20",X"B5",X"69",X"90",X"E2",X"20",X"9B",X"63",X"20",X"95",X"65",X"20",X"9B",X"63",X"4C",
		X"95",X"65",X"C9",X"00",X"F0",X"0C",X"98",X"10",X"06",X"20",X"8D",X"63",X"4C",X"C2",X"64",X"20",
		X"9B",X"63",X"20",X"95",X"65",X"A5",X"08",X"8D",X"64",X"18",X"A5",X"09",X"8D",X"65",X"18",X"A5",
		X"0A",X"8D",X"66",X"18",X"A5",X"0B",X"8D",X"67",X"18",X"8D",X"7E",X"18",X"20",X"B5",X"69",X"AD",
		X"18",X"18",X"90",X"05",X"C9",X"08",X"B0",X"06",X"60",X"C9",X"05",X"B0",X"01",X"60",X"A2",X"02",
		X"20",X"10",X"63",X"20",X"B5",X"69",X"90",X"08",X"06",X"1D",X"26",X"1E",X"06",X"19",X"26",X"1A",
		X"20",X"54",X"63",X"20",X"D6",X"68",X"B0",X"12",X"E6",X"A7",X"A5",X"2C",X"C5",X"BC",X"F0",X"01",
		X"60",X"20",X"54",X"63",X"20",X"D6",X"68",X"B0",X"01",X"60",X"24",X"CE",X"10",X"0B",X"09",X"00",
		X"30",X"0F",X"AD",X"2A",X"18",X"29",X"02",X"09",X"01",X"05",X"C5",X"85",X"C5",X"A9",X"30",X"85",
		X"C4",X"4C",X"BA",X"63",X"24",X"CE",X"10",X"39",X"A5",X"D1",X"C9",X"FF",X"F0",X"4B",X"AD",X"2A",
		X"18",X"4A",X"90",X"45",X"A5",X"B9",X"D0",X"41",X"A5",X"B8",X"38",X"E5",X"BA",X"F0",X"04",X"90",
		X"20",X"B0",X"36",X"A5",X"3A",X"29",X"07",X"D0",X"08",X"A9",X"01",X"05",X"C5",X"85",X"C5",X"D0",
		X"0B",X"A9",X"00",X"85",X"C5",X"20",X"10",X"68",X"49",X"40",X"85",X"BC",X"A9",X"40",X"85",X"C4",
		X"60",X"AD",X"2A",X"18",X"29",X"1F",X"24",X"3A",X"30",X"04",X"E5",X"BC",X"D0",X"02",X"65",X"BC",
		X"85",X"BC",X"A9",X"00",X"85",X"C5",X"4C",X"CB",X"63",X"20",X"10",X"68",X"85",X"BC",X"A9",X"80",
		X"85",X"C5",X"4C",X"CB",X"63",X"A5",X"D1",X"C9",X"20",X"B0",X"01",X"60",X"C9",X"FF",X"F0",X"16",
		X"A5",X"B9",X"D0",X"12",X"A5",X"B8",X"4A",X"D0",X"0D",X"A5",X"D0",X"C9",X"20",X"B0",X"EC",X"AD",
		X"E8",X"02",X"C9",X"24",X"B0",X"6D",X"20",X"10",X"68",X"A2",X"02",X"38",X"E5",X"2C",X"10",X"05",
		X"18",X"49",X"FF",X"69",X"02",X"C9",X"02",X"B0",X"5A",X"A5",X"26",X"D0",X"56",X"A5",X"12",X"D0",
		X"52",X"A9",X"7F",X"85",X"26",X"A9",X"05",X"85",X"BD",X"A5",X"15",X"29",X"F7",X"85",X"15",X"A5",
		X"2C",X"20",X"4B",X"5E",X"85",X"08",X"8A",X"85",X"B2",X"30",X"04",X"A9",X"00",X"F0",X"02",X"A9",
		X"FF",X"06",X"08",X"26",X"B2",X"2A",X"85",X"B3",X"A5",X"2C",X"20",X"4E",X"5E",X"85",X"08",X"8A",
		X"85",X"B6",X"30",X"04",X"A9",X"00",X"F0",X"02",X"A9",X"FF",X"06",X"08",X"26",X"B6",X"2A",X"85",
		X"B7",X"A5",X"2F",X"85",X"AA",X"A5",X"30",X"85",X"AB",X"A5",X"33",X"85",X"AE",X"A5",X"34",X"85",
		X"AF",X"A2",X"02",X"60",X"E6",X"A7",X"A9",X"00",X"CD",X"E4",X"02",X"A9",X"02",X"ED",X"E5",X"02",
		X"A9",X"00",X"2A",X"85",X"A6",X"25",X"CA",X"F0",X"03",X"4C",X"45",X"67",X"A5",X"2A",X"38",X"E5",
		X"BC",X"85",X"0A",X"10",X"05",X"18",X"49",X"FF",X"69",X"01",X"C9",X"40",X"B0",X"08",X"A2",X"02",
		X"24",X"0A",X"10",X"21",X"30",X"14",X"20",X"10",X"68",X"A2",X"02",X"85",X"0A",X"A5",X"BC",X"38",
		X"E5",X"0A",X"F0",X"15",X"10",X"0B",X"C9",X"FD",X"90",X"02",X"E6",X"BC",X"E6",X"BC",X"4C",X"79",
		X"66",X"C9",X"03",X"90",X"02",X"C6",X"BC",X"C6",X"BC",X"AD",X"EC",X"02",X"F0",X"24",X"A5",X"B9",
		X"D0",X"19",X"AD",X"00",X"0A",X"4A",X"4A",X"29",X"03",X"AA",X"BD",X"8A",X"38",X"18",X"F8",X"69",
		X"25",X"D8",X"38",X"E5",X"B8",X"30",X"04",X"C9",X"08",X"B0",X"02",X"A9",X"08",X"CD",X"E8",X"02",
		X"90",X"05",X"A5",X"BC",X"4C",X"BE",X"66",X"A5",X"C6",X"4A",X"4A",X"4A",X"4A",X"A5",X"C6",X"29",
		X"1F",X"85",X"08",X"A5",X"BC",X"B0",X"05",X"65",X"08",X"4C",X"BE",X"66",X"E5",X"08",X"85",X"2C",
		X"20",X"4E",X"5E",X"86",X"1D",X"48",X"A9",X"00",X"24",X"1D",X"10",X"02",X"A9",X"FF",X"85",X"1E",
		X"68",X"0A",X"26",X"1D",X"26",X"1E",X"0A",X"26",X"1D",X"26",X"1E",X"A5",X"2C",X"20",X"4B",X"5E",
		X"86",X"19",X"48",X"A9",X"00",X"24",X"19",X"10",X"02",X"A9",X"FF",X"85",X"1A",X"68",X"0A",X"26",
		X"19",X"26",X"1A",X"0A",X"26",X"19",X"26",X"1A",X"A5",X"2F",X"85",X"C0",X"A5",X"30",X"85",X"C1",
		X"A5",X"33",X"85",X"C2",X"A5",X"34",X"85",X"C3",X"A2",X"02",X"20",X"54",X"63",X"20",X"4E",X"5F",
		X"B0",X"1B",X"A2",X"02",X"20",X"D6",X"68",X"90",X"05",X"A6",X"A6",X"D0",X"11",X"60",X"A9",X"00",
		X"85",X"CA",X"AD",X"E4",X"02",X"0D",X"E5",X"02",X"F0",X"03",X"CE",X"E5",X"02",X"60",X"09",X"00",
		X"30",X"17",X"A5",X"C0",X"85",X"2F",X"A5",X"C1",X"85",X"30",X"A5",X"C2",X"85",X"33",X"A5",X"C3",
		X"85",X"34",X"E6",X"CA",X"60",X"EE",X"E5",X"02",X"60",X"A9",X"20",X"85",X"12",X"85",X"14",X"A9",
		X"02",X"85",X"C7",X"A9",X"FF",X"85",X"DF",X"A9",X"01",X"18",X"F8",X"65",X"BA",X"D8",X"85",X"BA",
		X"A2",X"00",X"8E",X"25",X"18",X"8E",X"27",X"18",X"20",X"99",X"61",X"A9",X"FF",X"85",X"0F",X"A5",
		X"15",X"29",X"FD",X"85",X"15",X"C6",X"CC",X"D0",X"02",X"E6",X"CD",X"60",X"A5",X"D4",X"F0",X"23",
		X"C9",X"30",X"90",X"05",X"A9",X"60",X"38",X"E5",X"D4",X"18",X"69",X"08",X"0A",X"0A",X"29",X"F0",
		X"8D",X"EA",X"02",X"C6",X"D4",X"C6",X"D4",X"D0",X"09",X"AD",X"2A",X"18",X"85",X"D3",X"A9",X"00",
		X"85",X"DE",X"60",X"A5",X"DE",X"F0",X"51",X"A5",X"D9",X"18",X"69",X"08",X"85",X"D9",X"A5",X"D3",
		X"F0",X"1D",X"18",X"A5",X"DA",X"65",X"D5",X"85",X"D5",X"A5",X"D6",X"65",X"DB",X"85",X"D6",X"A5",
		X"D7",X"18",X"65",X"DC",X"85",X"D7",X"A5",X"D8",X"65",X"DD",X"85",X"D8",X"C6",X"D3",X"60",X"AD",
		X"2A",X"18",X"85",X"DA",X"09",X"00",X"30",X"04",X"A9",X"00",X"F0",X"02",X"A9",X"FF",X"85",X"DB",
		X"AD",X"2A",X"18",X"85",X"DC",X"09",X"00",X"30",X"04",X"A9",X"00",X"F0",X"02",X"A9",X"FF",X"85",
		X"DD",X"AD",X"2A",X"18",X"4A",X"85",X"D3",X"60",X"A5",X"B8",X"4A",X"D0",X"01",X"60",X"A5",X"D3",
		X"D0",X"CA",X"AD",X"2A",X"18",X"85",X"D6",X"AD",X"2A",X"18",X"85",X"D8",X"E6",X"DE",X"D0",X"BF",
		X"A0",X"00",X"38",X"A5",X"2D",X"E5",X"2F",X"85",X"08",X"A5",X"2E",X"E5",X"30",X"85",X"09",X"10",
		X"04",X"20",X"49",X"61",X"C8",X"A5",X"08",X"85",X"0A",X"A5",X"09",X"85",X"0B",X"A5",X"09",X"38",
		X"A5",X"31",X"E5",X"33",X"85",X"08",X"A5",X"32",X"E5",X"34",X"85",X"09",X"10",X"0B",X"20",X"49",
		X"61",X"98",X"F0",X"03",X"C8",X"D0",X"02",X"A0",X"03",X"A5",X"08",X"C5",X"0A",X"D0",X"0D",X"A5",
		X"09",X"C5",X"0B",X"F0",X"03",X"38",X"B0",X"04",X"A9",X"20",X"D0",X"54",X"A5",X"09",X"E5",X"0B",
		X"08",X"90",X"1A",X"A5",X"08",X"8D",X"75",X"18",X"A5",X"09",X"8D",X"76",X"18",X"A5",X"0A",X"8D",
		X"6F",X"18",X"A5",X"0B",X"8D",X"70",X"18",X"8D",X"74",X"18",X"4C",X"94",X"68",X"A5",X"0A",X"8D",
		X"75",X"18",X"A5",X"0B",X"8D",X"76",X"18",X"A5",X"08",X"8D",X"6F",X"18",X"A5",X"09",X"8D",X"70",
		X"18",X"8D",X"74",X"18",X"20",X"80",X"5B",X"85",X"0C",X"AD",X"18",X"18",X"4A",X"66",X"0C",X"4A",
		X"66",X"0C",X"A6",X"0C",X"BD",X"85",X"37",X"28",X"90",X"06",X"85",X"0C",X"A9",X"40",X"E5",X"0C",
		X"AA",X"98",X"0A",X"A8",X"B9",X"BF",X"68",X"48",X"B9",X"BE",X"68",X"48",X"8A",X"60",X"D4",X"68",
		X"C5",X"68",X"CA",X"68",X"CF",X"68",X"18",X"49",X"FF",X"69",X"01",X"49",X"80",X"4C",X"D5",X"68",
		X"18",X"49",X"FF",X"69",X"01",X"60",X"18",X"86",X"08",X"B5",X"2D",X"8D",X"60",X"18",X"B5",X"2E",
		X"8D",X"61",X"18",X"B5",X"31",X"8D",X"62",X"18",X"B5",X"32",X"8D",X"63",X"18",X"A0",X"00",X"B9",
		X"CC",X"3F",X"30",X"67",X"B9",X"81",X"76",X"8D",X"64",X"18",X"B9",X"82",X"76",X"8D",X"65",X"18",
		X"B9",X"AB",X"76",X"8D",X"66",X"18",X"B9",X"AC",X"76",X"8D",X"7D",X"18",X"C1",X"00",X"AD",X"10",
		X"18",X"85",X"0C",X"AD",X"18",X"18",X"85",X"0D",X"8A",X"D0",X"08",X"A9",X"80",X"C5",X"0C",X"A9",
		X"04",X"D0",X"2E",X"B9",X"CC",X"3F",X"0A",X"AA",X"24",X"CB",X"10",X"1B",X"A5",X"0D",X"C9",X"80",
		X"6A",X"85",X"0B",X"A5",X"0C",X"6A",X"18",X"65",X"0C",X"85",X"0C",X"A5",X"0B",X"65",X"0D",X"85",
		X"0D",X"90",X"04",X"A6",X"08",X"B0",X"10",X"BD",X"95",X"69",X"C5",X"0C",X"BD",X"96",X"69",X"A6",
		X"08",X"E5",X"0D",X"A9",X"00",X"B0",X"3B",X"C8",X"C8",X"D0",X"94",X"A5",X"12",X"05",X"14",X"D0",
		X"31",X"8A",X"49",X"02",X"AA",X"B5",X"2D",X"8D",X"64",X"18",X"B5",X"2E",X"8D",X"65",X"18",X"B5",
		X"31",X"8D",X"66",X"18",X"B5",X"32",X"8D",X"7D",X"18",X"C1",X"00",X"AD",X"10",X"18",X"85",X"0C",
		X"AD",X"18",X"18",X"85",X"0D",X"A9",X"05",X"24",X"CB",X"10",X"02",X"A9",X"03",X"38",X"E5",X"0D",
		X"A9",X"FF",X"A6",X"08",X"60",X"40",X"03",X"40",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"C0",X"03",X"18",X"AD",X"EC",X"02",X"30",X"02",X"C9",X"05",X"60",X"A5",X"CD",
		X"D0",X"26",X"A5",X"B9",X"D0",X"0F",X"AD",X"00",X"0A",X"4A",X"4A",X"29",X"03",X"AA",X"A5",X"B8",
		X"DD",X"8A",X"38",X"90",X"13",X"AC",X"2A",X"18",X"98",X"4D",X"4A",X"03",X"8C",X"4A",X"03",X"4A",
		X"90",X"06",X"A9",X"02",X"85",X"D2",X"D0",X"3A",X"AD",X"2A",X"18",X"85",X"BC",X"A9",X"00",X"85",
		X"CB",X"85",X"14",X"A9",X"01",X"85",X"C4",X"85",X"D2",X"24",X"CE",X"10",X"20",X"A5",X"B9",X"D0",
		X"0D",X"38",X"A5",X"B8",X"E5",X"BA",X"90",X"15",X"F0",X"13",X"C9",X"07",X"90",X"02",X"A9",X"07",
		X"4A",X"F0",X"0A",X"AA",X"A9",X"0F",X"38",X"2A",X"CA",X"D0",X"FB",X"F0",X"28",X"A9",X"0F",X"4C",
		X"45",X"6A",X"EE",X"EC",X"02",X"A9",X"18",X"8D",X"E5",X"02",X"A9",X"00",X"8D",X"E4",X"02",X"A9",
		X"80",X"85",X"C5",X"A2",X"FF",X"8E",X"24",X"18",X"CA",X"8E",X"26",X"18",X"A9",X"FF",X"85",X"CB",
		X"AD",X"2A",X"18",X"29",X"0F",X"85",X"08",X"AD",X"2A",X"18",X"25",X"08",X"24",X"3A",X"70",X"02",
		X"49",X"FF",X"18",X"65",X"2A",X"85",X"08",X"20",X"4B",X"5E",X"85",X"0A",X"85",X"19",X"86",X"1A",
		X"8A",X"C9",X"80",X"6A",X"66",X"0A",X"C9",X"80",X"6A",X"66",X"0A",X"85",X"0B",X"A5",X"19",X"38",
		X"E5",X"0A",X"85",X"0A",X"A5",X"1A",X"E5",X"0B",X"AA",X"24",X"CB",X"30",X"0D",X"AD",X"2A",X"18",
		X"4A",X"08",X"8A",X"90",X"05",X"C9",X"80",X"6A",X"66",X"0A",X"85",X"0B",X"A5",X"08",X"20",X"4E",
		X"5E",X"85",X"08",X"85",X"1D",X"86",X"1E",X"8A",X"C9",X"80",X"6A",X"66",X"08",X"C9",X"80",X"6A",
		X"66",X"08",X"85",X"09",X"38",X"A5",X"1D",X"E5",X"08",X"85",X"08",X"A5",X"1E",X"E5",X"09",X"24",
		X"CB",X"30",X"08",X"28",X"90",X"05",X"C9",X"80",X"6A",X"66",X"08",X"85",X"09",X"18",X"A5",X"2D",
		X"65",X"0A",X"85",X"2F",X"A5",X"2E",X"65",X"0B",X"85",X"30",X"A5",X"31",X"18",X"65",X"08",X"85",
		X"33",X"A5",X"32",X"65",X"09",X"85",X"34",X"24",X"CB",X"10",X"07",X"20",X"10",X"68",X"85",X"2C",
		X"85",X"BC",X"A9",X"00",X"85",X"C9",X"85",X"D1",X"60",X"A2",X"3C",X"A9",X"35",X"20",X"5A",X"7A",
		X"A9",X"00",X"85",X"05",X"85",X"07",X"85",X"36",X"A9",X"0B",X"18",X"65",X"BF",X"85",X"BF",X"20",
		X"4E",X"5E",X"8A",X"C9",X"80",X"6A",X"85",X"04",X"85",X"35",X"10",X"06",X"A9",X"FF",X"85",X"05",
		X"85",X"36",X"A5",X"BF",X"20",X"4B",X"5E",X"8A",X"C9",X"80",X"6A",X"85",X"06",X"10",X"04",X"A9",
		X"FF",X"85",X"07",X"A9",X"A0",X"85",X"01",X"A9",X"3C",X"18",X"65",X"06",X"85",X"37",X"A9",X"01",
		X"65",X"07",X"85",X"38",X"20",X"AB",X"7A",X"A5",X"14",X"F0",X"09",X"A9",X"00",X"8D",X"25",X"18",
		X"8D",X"27",X"18",X"60",X"20",X"10",X"68",X"49",X"80",X"38",X"85",X"A6",X"A5",X"2A",X"E5",X"A6",
		X"85",X"A6",X"A5",X"BF",X"38",X"E5",X"A6",X"30",X"09",X"C9",X"0C",X"B0",X"05",X"A9",X"F0",X"8D",
		X"E9",X"02",X"A5",X"08",X"8D",X"64",X"18",X"A5",X"09",X"8D",X"65",X"18",X"A5",X"0A",X"8D",X"66",
		X"18",X"A5",X"0B",X"8D",X"67",X"18",X"8D",X"7E",X"18",X"C1",X"00",X"AD",X"10",X"18",X"85",X"0C",
		X"AD",X"18",X"18",X"8D",X"E8",X"02",X"AA",X"30",X"0B",X"4A",X"4A",X"4A",X"29",X"0F",X"49",X"AF",
		X"24",X"CB",X"30",X"02",X"A9",X"00",X"8D",X"25",X"18",X"8D",X"27",X"18",X"8A",X"8D",X"68",X"18",
		X"C9",X"80",X"90",X"1A",X"A9",X"00",X"85",X"C9",X"24",X"CB",X"10",X"0F",X"A5",X"D2",X"C9",X"04",
		X"90",X"06",X"20",X"E8",X"69",X"4C",X"5A",X"6C",X"20",X"22",X"6A",X"4C",X"5A",X"6C",X"AD",X"E9",
		X"02",X"D0",X"01",X"60",X"C9",X"F0",X"90",X"05",X"A9",X"01",X"20",X"85",X"79",X"A5",X"A6",X"20",
		X"4E",X"5E",X"8D",X"60",X"18",X"8E",X"61",X"18",X"A5",X"A6",X"20",X"4B",X"5E",X"8D",X"62",X"18",
		X"8E",X"63",X"18",X"A9",X"00",X"8D",X"64",X"18",X"A9",X"00",X"8D",X"65",X"18",X"A9",X"3C",X"8D",
		X"66",X"18",X"A9",X"01",X"8D",X"67",X"18",X"A9",X"00",X"8D",X"69",X"18",X"85",X"01",X"8D",X"6A",
		X"18",X"8D",X"71",X"18",X"20",X"80",X"5B",X"8D",X"77",X"18",X"AD",X"10",X"18",X"38",X"E5",X"35",
		X"85",X"04",X"AD",X"18",X"18",X"8D",X"79",X"18",X"E5",X"36",X"85",X"05",X"AD",X"10",X"18",X"38",
		X"E5",X"37",X"85",X"06",X"AD",X"18",X"18",X"E5",X"38",X"85",X"07",X"20",X"AB",X"7A",X"AD",X"E9",
		X"02",X"29",X"E0",X"20",X"8A",X"7A",X"A5",X"01",X"20",X"8A",X"7A",X"24",X"CE",X"30",X"05",X"2C",
		X"4B",X"03",X"30",X"0B",X"A9",X"02",X"25",X"C6",X"F0",X"05",X"A2",X"10",X"20",X"98",X"6C",X"A5",
		X"C9",X"D0",X"07",X"E6",X"C9",X"A9",X"10",X"20",X"85",X"79",X"AD",X"E9",X"02",X"F0",X"06",X"38",
		X"E9",X"08",X"8D",X"E9",X"02",X"60",X"A2",X"02",X"B5",X"24",X"F0",X"1E",X"30",X"1C",X"D6",X"24",
		X"18",X"B5",X"A8",X"75",X"B0",X"95",X"A8",X"B5",X"A9",X"75",X"B1",X"95",X"A9",X"B5",X"AC",X"18",
		X"75",X"B4",X"95",X"AC",X"B5",X"AD",X"75",X"B5",X"95",X"AD",X"CA",X"CA",X"F0",X"DA",X"60",X"6B",
		X"CB",X"6C",X"C0",X"6C",X"B5",X"6C",X"AA",X"6C",X"AD",X"00",X"0A",X"2A",X"2A",X"2A",X"2A",X"29",
		X"06",X"A8",X"B9",X"91",X"6C",X"48",X"B9",X"90",X"6C",X"48",X"60",X"BD",X"F6",X"70",X"85",X"3B",
		X"BD",X"F7",X"70",X"4C",X"D4",X"6C",X"BD",X"3A",X"6F",X"85",X"3B",X"BD",X"3B",X"6F",X"4C",X"D4",
		X"6C",X"BD",X"88",X"72",X"85",X"3B",X"BD",X"89",X"72",X"4C",X"D4",X"6C",X"BD",X"93",X"6D",X"85",
		X"3B",X"BD",X"94",X"6D",X"85",X"3C",X"A0",X"00",X"8A",X"C9",X"14",X"A9",X"02",X"90",X"02",X"A9",
		X"01",X"85",X"0D",X"B1",X"3B",X"C8",X"11",X"3B",X"F0",X"0E",X"20",X"6A",X"7A",X"A0",X"01",X"B1",
		X"3B",X"AA",X"88",X"B1",X"3B",X"20",X"8E",X"7A",X"A5",X"0D",X"20",X"81",X"7A",X"A0",X"02",X"A9",
		X"00",X"85",X"08",X"B1",X"3B",X"85",X"0A",X"29",X"7F",X"C8",X"84",X"0C",X"AA",X"BD",X"F0",X"33",
		X"A4",X"08",X"91",X"02",X"C8",X"BD",X"F1",X"33",X"91",X"02",X"C8",X"84",X"08",X"A4",X"0C",X"24",
		X"0A",X"10",X"E0",X"A4",X"08",X"88",X"20",X"76",X"7A",X"A9",X"01",X"4C",X"81",X"7A",X"20",X"6A",
		X"7A",X"A0",X"00",X"84",X"00",X"A2",X"5A",X"A9",X"20",X"20",X"8E",X"7A",X"A5",X"CC",X"F0",X"19",
		X"85",X"08",X"A0",X"00",X"AE",X"91",X"35",X"AD",X"90",X"35",X"91",X"02",X"8A",X"C8",X"91",X"02",
		X"C8",X"C6",X"08",X"D0",X"F2",X"88",X"20",X"76",X"7A",X"A2",X"18",X"20",X"98",X"6C",X"A0",X"00",
		X"A2",X"00",X"A9",X"D6",X"20",X"8E",X"7A",X"A9",X"B8",X"20",X"9E",X"7B",X"A2",X"0E",X"20",X"98",
		X"6C",X"A9",X"02",X"20",X"81",X"7A",X"A0",X"00",X"A2",X"00",X"A9",X"D6",X"20",X"8E",X"7A",X"AD",
		X"00",X"03",X"85",X"0A",X"AD",X"01",X"03",X"85",X"0B",X"A9",X"0A",X"20",X"9E",X"7B",X"A9",X"01",
		X"4C",X"81",X"7A",X"C3",X"6D",X"CE",X"6D",X"D4",X"6D",X"DB",X"6D",X"E1",X"6D",X"F6",X"6D",X"20",
		X"6E",X"40",X"6E",X"55",X"6E",X"65",X"6E",X"7F",X"6E",X"8A",X"6E",X"97",X"6E",X"A6",X"6E",X"B3",
		X"6E",X"B9",X"6E",X"C6",X"6E",X"D7",X"6E",X"E2",X"6E",X"ED",X"6E",X"FD",X"6E",X"0A",X"6F",X"1A",
		X"6F",X"2A",X"6F",X"92",X"4A",X"1E",X"30",X"1E",X"2E",X"46",X"00",X"3C",X"32",X"80",X"00",X"00",
		X"2C",X"1E",X"20",X"BC",X"00",X"00",X"38",X"26",X"22",X"24",X"BC",X"00",X"00",X"38",X"1E",X"16",
		X"B8",X"07",X"1A",X"1E",X"30",X"3C",X"1E",X"38",X"00",X"46",X"32",X"3E",X"38",X"00",X"26",X"30",
		X"26",X"3C",X"26",X"16",X"2C",X"BA",X"C4",X"10",X"1A",X"24",X"16",X"30",X"22",X"1E",X"00",X"2C",
		X"1E",X"3C",X"3C",X"1E",X"38",X"00",X"42",X"26",X"3C",X"24",X"00",X"38",X"26",X"22",X"24",X"3C",
		X"00",X"24",X"16",X"30",X"1C",X"00",X"1A",X"32",X"30",X"3C",X"38",X"32",X"2C",X"2C",X"1E",X"B8",
		X"D3",X"08",X"3A",X"1E",X"2C",X"1E",X"1A",X"3C",X"00",X"2C",X"1E",X"3C",X"3C",X"1E",X"38",X"00",
		X"42",X"26",X"3C",X"24",X"00",X"20",X"26",X"38",X"1E",X"00",X"18",X"3E",X"3C",X"3C",X"32",X"B0",
		X"20",X"46",X"24",X"26",X"22",X"24",X"00",X"3A",X"1A",X"32",X"38",X"1E",X"00",X"00",X"00",X"00",
		X"00",X"00",X"02",X"02",X"82",X"92",X"5A",X"1E",X"30",X"1E",X"2E",X"46",X"00",X"26",X"30",X"00",
		X"38",X"16",X"30",X"22",X"9E",X"92",X"52",X"2E",X"32",X"3C",X"26",X"32",X"30",X"00",X"18",X"2C",
		X"32",X"1A",X"2A",X"1E",X"1C",X"00",X"18",X"46",X"00",X"32",X"18",X"28",X"1E",X"1A",X"BC",X"E4",
		X"18",X"22",X"16",X"2E",X"1E",X"00",X"32",X"40",X"1E",X"B8",X"DE",X"00",X"34",X"38",X"1E",X"3A",
		X"3A",X"00",X"3A",X"3C",X"16",X"38",X"BC",X"20",X"50",X"3A",X"1A",X"32",X"38",X"1E",X"00",X"00",
		X"00",X"00",X"00",X"02",X"02",X"82",X"E4",X"28",X"24",X"26",X"22",X"24",X"00",X"3A",X"1A",X"32",
		X"38",X"1E",X"BA",X"00",X"00",X"02",X"02",X"02",X"80",X"C0",X"18",X"22",X"38",X"1E",X"16",X"3C",
		X"00",X"3A",X"1A",X"32",X"38",X"9E",X"CE",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"00",X"00",X"00",X"00",X"00",X"BA",X"CE",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"84",X"CE",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"3A",X"00",X"84",X"CE",X"00",X"00",
		X"00",X"1A",X"32",X"26",X"30",X"00",X"00",X"00",X"00",X"34",X"2C",X"16",X"C6",X"DC",X"EA",X"26",
		X"30",X"3A",X"1E",X"38",X"3C",X"00",X"1A",X"32",X"26",X"B0",X"A9",X"BA",X"18",X"32",X"30",X"3E",
		X"3A",X"00",X"3C",X"16",X"30",X"2A",X"00",X"16",X"3C",X"80",X"00",X"00",X"02",X"02",X"02",X"00",
		X"16",X"30",X"1C",X"00",X"04",X"02",X"02",X"02",X"02",X"82",X"D6",X"C4",X"4E",X"50",X"00",X"00",
		X"16",X"3C",X"16",X"38",X"26",X"00",X"04",X"14",X"12",X"82",X"6A",X"6F",X"73",X"6F",X"7D",X"6F",
		X"87",X"6F",X"91",X"6F",X"A9",X"6F",X"DF",X"6F",X"09",X"70",X"22",X"70",X"33",X"70",X"47",X"70",
		X"56",X"70",X"97",X"6E",X"69",X"70",X"B3",X"6E",X"7A",X"70",X"87",X"70",X"9B",X"70",X"A7",X"70",
		X"B3",X"70",X"C6",X"70",X"DD",X"70",X"E7",X"70",X"2A",X"6F",X"88",X"4A",X"1E",X"30",X"30",X"1E",
		X"2E",X"26",X"80",X"00",X"00",X"16",X"00",X"22",X"16",X"3E",X"1A",X"24",X"9E",X"00",X"00",X"16",
		X"00",X"1C",X"38",X"32",X"26",X"3C",X"9E",X"00",X"00",X"1C",X"1E",X"38",X"38",X"26",X"1E",X"38",
		X"9E",X"07",X"1A",X"1A",X"32",X"2E",X"34",X"32",X"3A",X"1E",X"38",X"00",X"40",X"32",X"3A",X"00",
		X"26",X"30",X"26",X"3C",X"26",X"16",X"2C",X"1E",X"BA",X"B4",X"10",X"1A",X"24",X"32",X"26",X"3A",
		X"26",X"3A",X"3A",X"1E",X"48",X"00",X"40",X"32",X"3C",X"38",X"1E",X"00",X"2C",X"1E",X"3C",X"3C",
		X"38",X"1E",X"00",X"16",X"40",X"1E",X"1A",X"00",X"2C",X"1E",X"00",X"1A",X"32",X"30",X"3C",X"38",
		X"32",X"2C",X"1E",X"3E",X"38",X"00",X"1C",X"1E",X"00",X"1C",X"38",X"32",X"26",X"3C",X"9E",X"BF",
		X"08",X"16",X"34",X"34",X"3E",X"46",X"1E",X"38",X"00",X"3A",X"3E",X"38",X"00",X"20",X"1E",X"3E",
		X"00",X"34",X"32",X"3E",X"38",X"00",X"3A",X"1E",X"2C",X"1E",X"1A",X"3C",X"26",X"32",X"30",X"00",
		X"1C",X"1E",X"00",X"2C",X"1E",X"3C",X"3C",X"38",X"9E",X"20",X"46",X"2E",X"1E",X"26",X"2C",X"2C",
		X"1E",X"3E",X"38",X"00",X"3A",X"1A",X"32",X"38",X"1E",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"02",X"82",X"88",X"5A",X"1E",X"30",X"30",X"1E",X"2E",X"26",X"00",X"16",X"00",X"34",X"32",X"38",
		X"3C",X"1E",X"9E",X"88",X"52",X"16",X"3C",X"3C",X"1E",X"30",X"3C",X"26",X"32",X"30",X"00",X"32",
		X"18",X"3A",X"3C",X"16",X"1A",X"2C",X"9E",X"E0",X"18",X"20",X"26",X"30",X"00",X"1C",X"1E",X"00",
		X"34",X"16",X"38",X"3C",X"26",X"9E",X"CE",X"00",X"16",X"34",X"34",X"3E",X"46",X"1E",X"48",X"00",
		X"3A",X"3E",X"38",X"00",X"3A",X"3C",X"16",X"38",X"BC",X"DC",X"28",X"2E",X"1E",X"26",X"2C",X"2C",
		X"1E",X"3E",X"38",X"3A",X"00",X"3A",X"1A",X"32",X"38",X"9E",X"C0",X"18",X"3A",X"1A",X"32",X"38",
		X"1E",X"00",X"1E",X"2C",X"1E",X"40",X"9E",X"C6",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BA",X"C6",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"84",X"C6",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3A",X"00",X"84",X"C6",X"00",X"00",X"00",X"34",X"26",X"1E",X"1A",X"1E",X"00",X"00",X"00",X"00",
		X"28",X"32",X"3E",X"1E",X"3E",X"B8",X"CA",X"EA",X"26",X"30",X"3C",X"38",X"32",X"1C",X"3E",X"26",
		X"38",X"1E",X"00",X"2C",X"1E",X"3A",X"00",X"34",X"26",X"1E",X"1A",X"1E",X"BA",X"BE",X"BA",X"18",
		X"32",X"30",X"3E",X"3A",X"00",X"16",X"80",X"00",X"00",X"02",X"02",X"02",X"00",X"1E",X"3C",X"00",
		X"04",X"02",X"02",X"02",X"02",X"82",X"26",X"71",X"34",X"71",X"44",X"71",X"52",X"71",X"59",X"71",
		X"6E",X"71",X"94",X"71",X"B5",X"71",X"CD",X"71",X"DF",X"71",X"00",X"72",X"11",X"72",X"1F",X"72",
		X"2F",X"72",X"B3",X"6E",X"38",X"72",X"87",X"70",X"9B",X"70",X"A7",X"70",X"48",X"72",X"5B",X"72",
		X"6B",X"72",X"7A",X"72",X"2A",X"6F",X"85",X"4A",X"1E",X"30",X"1E",X"2E",X"26",X"22",X"32",X"00",
		X"2E",X"3E",X"46",X"80",X"00",X"00",X"16",X"00",X"2C",X"16",X"00",X"26",X"48",X"36",X"3E",X"26",
		X"1E",X"38",X"1C",X"96",X"00",X"00",X"16",X"00",X"2C",X"16",X"00",X"1C",X"1E",X"38",X"1E",X"1A",
		X"24",X"96",X"00",X"00",X"16",X"3C",X"38",X"16",X"BA",X"02",X"1A",X"22",X"38",X"16",X"18",X"1E",
		X"00",X"3A",X"3E",X"3A",X"00",X"26",X"30",X"26",X"1A",X"26",X"16",X"2C",X"1E",X"BA",X"C2",X"10",
		X"3A",X"1E",X"2C",X"1E",X"1A",X"1A",X"26",X"32",X"30",X"1E",X"00",X"2C",X"1E",X"3C",X"38",X"16",
		X"00",X"1A",X"32",X"30",X"00",X"1A",X"32",X"30",X"3C",X"38",X"32",X"2C",X"00",X"1C",X"1E",X"38",
		X"1E",X"1A",X"24",X"B2",X"C9",X"08",X"22",X"38",X"16",X"18",X"1E",X"2C",X"16",X"00",X"1A",X"32",
		X"30",X"00",X"1E",X"2C",X"00",X"18",X"32",X"3C",X"32",X"30",X"00",X"1C",X"1E",X"00",X"1C",X"26",
		X"3A",X"34",X"16",X"38",X"B2",X"20",X"46",X"34",X"3E",X"30",X"3C",X"32",X"3A",X"00",X"2E",X"16",
		X"46",X"32",X"38",X"1E",X"3A",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"82",X"85",X"5A",X"1E",
		X"30",X"1E",X"2E",X"26",X"22",X"32",X"00",X"1E",X"30",X"00",X"38",X"16",X"30",X"22",X"B2",X"85",
		X"52",X"2E",X"32",X"40",X"26",X"2E",X"26",X"1E",X"30",X"3C",X"32",X"00",X"18",X"2C",X"32",X"36",
		X"3E",X"1E",X"16",X"1C",X"32",X"00",X"34",X"32",X"38",X"00",X"32",X"18",X"28",X"1E",X"3C",X"B2",
		X"D8",X"18",X"28",X"3E",X"1E",X"22",X"32",X"00",X"3C",X"1E",X"38",X"2E",X"26",X"30",X"16",X"1C",
		X"B2",X"DE",X"00",X"34",X"3E",X"2C",X"3A",X"16",X"38",X"00",X"3A",X"3C",X"16",X"38",X"BC",X"20",
		X"50",X"34",X"3E",X"30",X"3C",X"32",X"3A",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"82",X"F2",
		X"28",X"38",X"1E",X"1A",X"32",X"38",X"1C",X"BA",X"A8",X"18",X"34",X"3E",X"30",X"3C",X"32",X"3A",
		X"00",X"22",X"38",X"16",X"30",X"1C",X"1E",X"BA",X"C6",X"00",X"00",X"00",X"20",X"26",X"1A",X"24",
		X"16",X"00",X"00",X"00",X"00",X"00",X"28",X"1E",X"3E",X"22",X"B2",X"D8",X"EA",X"26",X"30",X"3A",
		X"1E",X"38",X"3C",X"1E",X"00",X"20",X"26",X"1A",X"24",X"16",X"BA",X"B2",X"BA",X"40",X"26",X"1C",
		X"16",X"00",X"1E",X"44",X"3C",X"38",X"16",X"00",X"16",X"80",X"00",X"00",X"02",X"02",X"02",X"00",
		X"46",X"00",X"04",X"02",X"02",X"02",X"02",X"82",X"B8",X"72",X"C5",X"72",X"CC",X"72",X"D4",X"72",
		X"DC",X"72",X"FA",X"72",X"32",X"73",X"63",X"73",X"7D",X"73",X"95",X"73",X"A9",X"73",X"B4",X"73",
		X"C9",X"73",X"DB",X"73",X"B3",X"6E",X"EE",X"73",X"05",X"74",X"19",X"74",X"26",X"74",X"33",X"74",
		X"46",X"74",X"56",X"74",X"62",X"74",X"2A",X"6F",X"85",X"4A",X"22",X"1E",X"22",X"30",X"1E",X"38",
		X"00",X"40",X"32",X"30",X"80",X"00",X"00",X"2C",X"26",X"30",X"2A",X"BA",X"00",X"00",X"38",X"1E",
		X"1A",X"24",X"3C",X"BA",X"00",X"00",X"24",X"26",X"30",X"3C",X"1E",X"B0",X"20",X"1A",X"22",X"1E",
		X"18",X"1E",X"30",X"00",X"3A",X"26",X"1E",X"00",X"26",X"24",X"38",X"1E",X"00",X"26",X"30",X"26",
		X"3C",X"26",X"16",X"2C",X"1E",X"30",X"00",X"1E",X"26",X"B0",X"B2",X"10",X"42",X"16",X"1E",X"24",
		X"2C",X"1E",X"30",X"00",X"3A",X"26",X"1E",X"00",X"1C",X"1E",X"30",X"00",X"18",X"3E",X"1A",X"24",
		X"3A",X"3C",X"16",X"18",X"1E",X"30",X"00",X"2E",X"26",X"3C",X"00",X"1C",X"1E",X"2E",X"00",X"38",
		X"1E",X"1A",X"24",X"3C",X"1E",X"30",X"00",X"3A",X"3C",X"1E",X"3E",X"1E",X"38",X"22",X"38",X"26",
		X"20",X"A0",X"C4",X"08",X"22",X"1E",X"18",X"1E",X"30",X"00",X"3A",X"26",X"1E",X"00",X"1C",X"1E",
		X"30",X"00",X"18",X"3E",X"1A",X"24",X"3A",X"3C",X"16",X"18",X"1E",X"30",X"00",X"2E",X"26",X"3C",
		X"00",X"1C",X"1E",X"2E",X"00",X"20",X"1E",X"3E",X"1E",X"38",X"2A",X"30",X"32",X"34",X"20",X"00",
		X"1E",X"26",X"B0",X"20",X"46",X"18",X"1E",X"3A",X"3C",X"1E",X"00",X"34",X"3E",X"30",X"2A",X"3C",
		X"48",X"16",X"24",X"2C",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"82",X"85",X"5A",X"22",
		X"1E",X"22",X"30",X"1E",X"38",X"00",X"26",X"2E",X"00",X"20",X"1E",X"3E",X"1E",X"38",X"18",X"1E",
		X"38",X"1E",X"26",X"1A",X"A4",X"85",X"52",X"18",X"1E",X"42",X"1E",X"22",X"3E",X"30",X"22",X"00",
		X"18",X"2C",X"32",X"1A",X"2A",X"26",X"1E",X"38",X"BC",X"E4",X"18",X"3A",X"34",X"26",X"1E",X"2C",
		X"1E",X"30",X"1C",X"9E",X"C6",X"00",X"3A",X"3C",X"16",X"38",X"3C",X"2A",X"30",X"32",X"34",X"20",
		X"00",X"1C",X"38",X"3E",X"1E",X"1A",X"2A",X"1E",X"B0",X"20",X"50",X"34",X"3E",X"30",X"2A",X"3C",
		X"48",X"16",X"24",X"2C",X"00",X"00",X"00",X"00",X"02",X"02",X"82",X"D6",X"28",X"24",X"32",X"1E",
		X"1A",X"24",X"3A",X"3C",X"1E",X"38",X"22",X"1E",X"18",X"30",X"26",X"3A",X"3A",X"9E",X"98",X"18",
		X"22",X"38",X"32",X"3A",X"3A",X"16",X"38",X"3C",X"26",X"22",X"1E",X"3A",X"00",X"1E",X"38",X"22",
		X"1E",X"18",X"30",X"26",X"BA",X"CA",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"9E",X"CA",X"00",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"84",X"CA",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"00",X"84",X"CA",X"00",X"00",X"00",X"2E",X"3E",X"1E",X"30",X"48",X"1E",X"00",X"00",X"00",
		X"00",X"3A",X"34",X"26",X"1E",X"AC",X"D8",X"EA",X"22",X"1E",X"2C",X"1C",X"00",X"1E",X"26",X"30",
		X"42",X"1E",X"38",X"20",X"1E",X"B0",X"B7",X"BA",X"18",X"32",X"30",X"3E",X"3A",X"00",X"18",X"1E",
		X"26",X"80",X"00",X"00",X"02",X"02",X"02",X"00",X"3E",X"30",X"1C",X"00",X"04",X"02",X"02",X"02",
		X"02",X"82",X"CB",X"74",X"D7",X"74",X"E9",X"74",X"19",X"75",X"25",X"75",X"25",X"75",X"25",X"75",
		X"25",X"75",X"25",X"75",X"25",X"75",X"25",X"75",X"25",X"75",X"CB",X"74",X"2D",X"75",X"3B",X"75",
		X"D7",X"74",X"5C",X"75",X"6A",X"75",X"3E",X"75",X"2D",X"75",X"6A",X"75",X"5C",X"75",X"7C",X"75",
		X"2F",X"76",X"6A",X"75",X"E6",X"75",X"5C",X"75",X"DC",X"75",X"5C",X"75",X"E6",X"75",X"49",X"76",
		X"61",X"76",X"B5",X"75",X"FF",X"75",X"00",X"00",X"00",X"00",X"F4",X"75",X"F4",X"75",X"F4",X"75",
		X"F4",X"75",X"F4",X"75",X"F4",X"75",X"F4",X"75",X"F4",X"75",X"DD",X"03",X"A1",X"24",X"0C",X"04",
		X"1C",X"24",X"14",X"1C",X"12",X"0C",X"FF",X"03",X"A1",X"0C",X"14",X"1C",X"04",X"24",X"2C",X"34",
		X"3C",X"24",X"2A",X"0C",X"12",X"34",X"3A",X"1C",X"FF",X"BB",X"A1",X"B4",X"62",X"6C",X"72",X"A4",
		X"94",X"7C",X"74",X"8C",X"84",X"9C",X"AC",X"8C",X"7A",X"84",X"9A",X"94",X"A2",X"AC",X"1B",X"04",
		X"24",X"3C",X"34",X"14",X"1C",X"3C",X"5C",X"54",X"34",X"2C",X"4C",X"54",X"6C",X"4C",X"44",X"5C",
		X"64",X"44",X"24",X"2C",X"0C",X"14",X"0A",X"04",X"FF",X"03",X"E1",X"24",X"0C",X"04",X"1C",X"24",
		X"14",X"1C",X"12",X"0C",X"FF",X"03",X"81",X"0C",X"12",X"1C",X"22",X"2C",X"FF",X"03",X"A1",X"0C",
		X"14",X"1C",X"04",X"24",X"2C",X"34",X"3C",X"24",X"3A",X"1C",X"FF",X"03",X"05",X"FF",X"03",X"A1",
		X"0C",X"14",X"1C",X"04",X"24",X"2C",X"0C",X"2A",X"14",X"1A",X"24",X"32",X"64",X"54",X"3C",X"34",
		X"4C",X"44",X"5C",X"6C",X"4C",X"3A",X"44",X"5A",X"54",X"62",X"6C",X"FF",X"03",X"A1",X"1C",X"2C",
		X"14",X"04",X"0C",X"14",X"2C",X"24",X"0C",X"22",X"1C",X"FF",X"03",X"A1",X"0C",X"14",X"1C",X"04",
		X"24",X"34",X"3C",X"2C",X"24",X"2A",X"0C",X"3A",X"14",X"1A",X"34",X"FF",X"6B",X"A1",X"64",X"34",
		X"04",X"0C",X"3C",X"44",X"4C",X"54",X"5C",X"34",X"3C",X"64",X"44",X"14",X"1C",X"4C",X"64",X"54",
		X"24",X"2C",X"5C",X"64",X"C3",X"E1",X"BC",X"B4",X"C4",X"CC",X"BC",X"CA",X"B4",X"0A",X"A1",X"14",
		X"1A",X"24",X"2A",X"04",X"93",X"9C",X"A4",X"AC",X"94",X"74",X"7C",X"84",X"8C",X"74",X"7A",X"9C",
		X"A2",X"84",X"8A",X"AC",X"FF",X"83",X"A1",X"44",X"4C",X"84",X"54",X"5C",X"84",X"64",X"6C",X"84",
		X"74",X"7C",X"84",X"03",X"3C",X"7C",X"44",X"04",X"0C",X"4C",X"54",X"14",X"1C",X"5C",X"64",X"24",
		X"2C",X"6C",X"74",X"34",X"3C",X"32",X"2C",X"22",X"1C",X"12",X"0C",X"FF",X"03",X"A1",X"14",X"0C",
		X"1C",X"04",X"0C",X"12",X"1C",X"FF",X"0B",X"A1",X"14",X"1C",X"3C",X"34",X"2C",X"24",X"04",X"0C",
		X"2C",X"32",X"14",X"FF",X"3B",X"A1",X"00",X"08",X"10",X"18",X"20",X"28",X"30",X"38",X"FF",X"03",
		X"A1",X"0C",X"24",X"04",X"1C",X"14",X"2C",X"1C",X"12",X"0C",X"22",X"2C",X"4B",X"54",X"34",X"74",
		X"6C",X"4C",X"44",X"3C",X"34",X"5C",X"64",X"44",X"62",X"6C",X"72",X"5C",X"9B",X"B4",X"AC",X"A4",
		X"84",X"7C",X"94",X"8C",X"84",X"7A",X"9C",X"B2",X"94",X"8A",X"AC",X"BA",X"E1",X"C4",X"FF",X"03",
		X"F1",X"0C",X"14",X"1C",X"24",X"2C",X"34",X"04",X"3A",X"44",X"4C",X"54",X"5C",X"3C",X"62",X"6C",
		X"74",X"7C",X"64",X"82",X"8C",X"94",X"9C",X"84",X"FF",X"03",X"0C",X"14",X"1C",X"24",X"2C",X"34",
		X"3C",X"44",X"4C",X"54",X"5C",X"64",X"6C",X"74",X"7C",X"3C",X"84",X"8C",X"94",X"9C",X"A4",X"04",
		X"FF",X"0B",X"04",X"2C",X"24",X"1C",X"14",X"0C",X"1C",X"3C",X"34",X"0C",X"4A",X"44",X"5C",X"54",
		X"4C",X"72",X"B4",X"BC",X"C4",X"64",X"6C",X"74",X"7C",X"84",X"8C",X"94",X"9C",X"A4",X"AC",X"B4",
		X"FF",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"80",X"00",X"80",X"00",X"80",X"00",
		X"40",X"00",X"30",X"00",X"C0",X"00",X"F7",X"00",X"C8",X"00",X"D8",X"00",X"94",X"00",X"98",X"00",
		X"E8",X"00",X"70",X"00",X"78",X"00",X"40",X"00",X"24",X"00",X"2C",X"00",X"20",X"00",X"40",X"00",
		X"80",X"00",X"80",X"00",X"80",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"18",X"00",
		X"44",X"00",X"40",X"00",X"8C",X"00",X"0C",X"00",X"E8",X"00",X"E4",X"00",X"9C",X"00",X"CC",X"00",
		X"B4",X"00",X"BC",X"00",X"F4",X"79",X"E0",X"00",X"00",X"14",X"20",X"00",X"E0",X"00",X"00",X"0F",
		X"20",X"00",X"A0",X"02",X"80",X"0C",X"58",X"00",X"60",X"04",X"C0",X"0D",X"90",X"00",X"40",X"06",
		X"80",X"0C",X"C8",X"00",X"00",X"08",X"00",X"0F",X"00",X"01",X"00",X"08",X"00",X"14",X"00",X"01",
		X"A0",X"02",X"80",X"11",X"58",X"00",X"A0",X"02",X"40",X"10",X"58",X"00",X"60",X"04",X"80",X"11",
		X"90",X"00",X"40",X"06",X"40",X"10",X"C8",X"00",X"40",X"06",X"80",X"11",X"C8",X"00",X"E0",X"00",
		X"80",X"0C",X"20",X"00",X"20",X"00",X"C0",X"08",X"58",X"00",X"E0",X"00",X"00",X"05",X"20",X"00",
		X"00",X"08",X"C0",X"08",X"00",X"01",X"80",X"03",X"00",X"0A",X"70",X"00",X"00",X"04",X"C0",X"08",
		X"80",X"00",X"80",X"03",X"80",X"07",X"70",X"00",X"40",X"05",X"C0",X"08",X"A8",X"00",X"7F",X"E0",
		X"00",X"80",X"02",X"20",X"00",X"40",X"06",X"40",X"01",X"C8",X"00",X"40",X"06",X"80",X"FD",X"C8",
		X"00",X"E0",X"00",X"40",X"FC",X"20",X"00",X"40",X"06",X"00",X"FB",X"C8",X"00",X"40",X"06",X"40",
		X"F7",X"C8",X"00",X"E0",X"00",X"40",X"F7",X"20",X"00",X"E0",X"00",X"00",X"F1",X"20",X"00",X"C0",
		X"01",X"C0",X"EA",X"38",X"00",X"A0",X"02",X"80",X"EE",X"58",X"00",X"80",X"03",X"80",X"EE",X"70",
		X"00",X"60",X"04",X"00",X"EC",X"90",X"00",X"40",X"05",X"80",X"EE",X"A8",X"00",X"40",X"06",X"80",
		X"EE",X"C8",X"00",X"20",X"07",X"C0",X"EA",X"E0",X"00",X"00",X"08",X"00",X"F1",X"00",X"01",X"A0",
		X"02",X"C0",X"F4",X"58",X"00",X"00",X"08",X"C0",X"F4",X"00",X"01",X"00",X"08",X"80",X"07",X"00",
		X"01",X"40",X"06",X"80",X"07",X"C8",X"00",X"40",X"06",X"C0",X"03",X"C8",X"00",X"97",X"00",X"F8",
		X"C0",X"12",X"00",X"FF",X"00",X"F8",X"C0",X"08",X"00",X"FF",X"C0",X"F9",X"C0",X"0D",X"38",X"FF",
		X"20",X"FF",X"C0",X"08",X"E0",X"FF",X"20",X"FF",X"C0",X"12",X"E0",X"FF",X"60",X"FD",X"C0",X"0D",
		X"A8",X"FF",X"00",X"F8",X"40",X"01",X"00",X"FF",X"20",X"FF",X"40",X"01",X"E0",X"FF",X"C0",X"F9",
		X"40",X"06",X"38",X"FF",X"C0",X"F9",X"C0",X"03",X"38",X"FF",X"60",X"FD",X"C0",X"03",X"A8",X"FF",
		X"60",X"FD",X"40",X"06",X"A8",X"FF",X"00",X"F8",X"00",X"00",X"00",X"FF",X"A0",X"FB",X"80",X"FD",
		X"70",X"FF",X"00",X"F8",X"00",X"F6",X"00",X"FF",X"E0",X"F8",X"C0",X"EF",X"20",X"FF",X"C0",X"F9",
		X"80",X"F3",X"38",X"FF",X"C0",X"FA",X"80",X"F3",X"58",X"FF",X"A0",X"FB",X"00",X"F1",X"70",X"FF",
		X"80",X"FC",X"80",X"F3",X"90",X"FF",X"60",X"FD",X"80",X"F3",X"A8",X"FF",X"40",X"FE",X"C0",X"EF",
		X"C8",X"FF",X"20",X"FF",X"00",X"F6",X"E0",X"FF",X"A0",X"FB",X"80",X"F8",X"70",X"FF",X"20",X"FF",
		X"00",X"00",X"E0",X"FF",X"00",X"00",X"15",X"1B",X"2D",X"57",X"00",X"00",X"21",X"27",X"00",X"00",
		X"00",X"00",X"61",X"67",X"00",X"00",X"01",X"0F",X"85",X"8F",X"00",X"00",X"95",X"A7",X"00",X"00",
		X"AD",X"D3",X"D9",X"D3",X"00",X"00",X"00",X"40",X"02",X"FF",X"18",X"40",X"02",X"FF",X"18",X"40",
		X"02",X"FF",X"18",X"00",X"00",X"A3",X"30",X"00",X"03",X"00",X"00",X"23",X"10",X"00",X"01",X"00",
		X"00",X"A3",X"10",X"00",X"01",X"00",X"00",X"10",X"01",X"00",X"20",X"00",X"00",X"C1",X"10",X"FF",
		X"02",X"00",X"00",X"C0",X"01",X"F6",X"06",X"84",X"01",X"09",X"0C",X"F0",X"01",X"F8",X"0C",X"90",
		X"01",X"07",X"0C",X"E4",X"01",X"FA",X"0C",X"9C",X"01",X"05",X"0C",X"D8",X"01",X"FC",X"0C",X"A8",
		X"01",X"03",X"0C",X"CC",X"01",X"FE",X"0C",X"B4",X"01",X"01",X"0C",X"00",X"00",X"AB",X"04",X"FF",
		X"09",X"A2",X"27",X"FF",X"02",X"00",X"00",X"10",X"70",X"00",X"02",X"00",X"00",X"A2",X"20",X"00",
		X"01",X"A0",X"20",X"00",X"01",X"A2",X"20",X"00",X"01",X"A0",X"20",X"00",X"01",X"A2",X"20",X"00",
		X"01",X"A0",X"20",X"00",X"01",X"A2",X"20",X"00",X"01",X"00",X"00",X"30",X"01",X"FC",X"0C",X"30",
		X"01",X"FC",X"0C",X"00",X"00",X"A3",X"02",X"00",X"0C",X"00",X"00",X"40",X"01",X"FE",X"10",X"20",
		X"01",X"02",X"10",X"40",X"01",X"FE",X"10",X"20",X"01",X"02",X"10",X"00",X"00",X"A1",X"10",X"00",
		X"04",X"00",X"00",X"D9",X"30",X"00",X"01",X"A2",X"30",X"00",X"01",X"90",X"30",X"00",X"01",X"80",
		X"30",X"00",X"01",X"90",X"30",X"00",X"01",X"A2",X"30",X"00",X"01",X"90",X"30",X"00",X"01",X"80",
		X"30",X"00",X"02",X"A2",X"30",X"00",X"04",X"00",X"00",X"A7",X"30",X"00",X"0D",X"00",X"00",X"6C",
		X"30",X"00",X"01",X"51",X"30",X"00",X"01",X"48",X"30",X"00",X"01",X"40",X"30",X"00",X"01",X"48",
		X"30",X"00",X"01",X"51",X"30",X"00",X"01",X"48",X"30",X"00",X"01",X"40",X"30",X"00",X"02",X"51",
		X"30",X"00",X"04",X"00",X"00",X"48",X"8A",X"48",X"98",X"48",X"BA",X"BD",X"03",X"01",X"F0",X"06",
		X"A2",X"08",X"0A",X"CA",X"90",X"FC",X"8A",X"0A",X"0A",X"69",X"03",X"A8",X"C0",X"27",X"B0",X"13",
		X"A2",X"03",X"B9",X"64",X"78",X"F0",X"08",X"95",X"EF",X"A9",X"01",X"95",X"F7",X"95",X"FB",X"88",
		X"CA",X"10",X"EF",X"68",X"A8",X"68",X"AA",X"68",X"60",X"A2",X"03",X"B5",X"F7",X"F0",X"1D",X"D6",
		X"F7",X"D0",X"47",X"B4",X"EF",X"F0",X"43",X"D6",X"FB",X"D0",X"32",X"B9",X"86",X"78",X"95",X"F3",
		X"B9",X"87",X"78",X"95",X"F7",X"D0",X"17",X"95",X"EF",X"8A",X"D0",X"2E",X"AD",X"85",X"78",X"95",
		X"F3",X"9D",X"20",X"18",X"A9",X"00",X"95",X"EF",X"CA",X"10",X"D0",X"4C",X"18",X"7A",X"B9",X"89",
		X"78",X"95",X"FB",X"B5",X"EF",X"18",X"69",X"04",X"95",X"EF",X"4C",X"0A",X"7A",X"B9",X"83",X"78",
		X"95",X"F7",X"B5",X"F3",X"18",X"79",X"84",X"78",X"95",X"F3",X"B5",X"F3",X"9D",X"20",X"18",X"AD",
		X"84",X"78",X"8D",X"28",X"18",X"CA",X"10",X"A3",X"60",X"A9",X"C0",X"D0",X"05",X"20",X"6A",X"7A",
		X"A9",X"20",X"A0",X"00",X"91",X"02",X"4C",X"C7",X"7A",X"90",X"04",X"29",X"0F",X"F0",X"05",X"29",
		X"0F",X"18",X"69",X"01",X"08",X"0A",X"A0",X"00",X"AA",X"BD",X"F0",X"33",X"91",X"02",X"BD",X"F1",
		X"33",X"C8",X"91",X"02",X"20",X"76",X"7A",X"28",X"60",X"4A",X"29",X"0F",X"09",X"E0",X"A0",X"01",
		X"91",X"02",X"88",X"8A",X"6A",X"91",X"02",X"C8",X"D0",X"1C",X"4A",X"29",X"0F",X"09",X"A0",X"D0",
		X"ED",X"A4",X"01",X"09",X"60",X"AA",X"98",X"4C",X"6E",X"7A",X"A9",X"40",X"A2",X"80",X"A0",X"00",
		X"91",X"02",X"C8",X"8A",X"91",X"02",X"98",X"38",X"65",X"02",X"85",X"02",X"90",X"02",X"E6",X"03",
		X"60",X"A0",X"00",X"09",X"70",X"AA",X"98",X"4C",X"6E",X"7A",X"A8",X"A9",X"00",X"AA",X"84",X"01",
		X"A0",X"00",X"0A",X"90",X"01",X"88",X"84",X"05",X"0A",X"26",X"05",X"85",X"04",X"8A",X"0A",X"A0",
		X"00",X"90",X"01",X"88",X"84",X"07",X"0A",X"26",X"07",X"85",X"06",X"A2",X"04",X"A0",X"00",X"B5",
		X"02",X"91",X"02",X"B5",X"03",X"29",X"1F",X"C8",X"91",X"02",X"B5",X"00",X"C8",X"91",X"02",X"B5",
		X"01",X"45",X"01",X"29",X"1F",X"45",X"01",X"C8",X"91",X"02",X"D0",X"AA",X"A2",X"7F",X"9A",X"A9",
		X"00",X"8D",X"2F",X"18",X"D8",X"AA",X"95",X"00",X"E8",X"D0",X"FB",X"A0",X"07",X"8C",X"2F",X"18",
		X"9D",X"00",X"01",X"9D",X"00",X"02",X"9D",X"00",X"03",X"9D",X"00",X"20",X"9D",X"00",X"21",X"9D",
		X"00",X"22",X"9D",X"00",X"23",X"9D",X"00",X"24",X"9D",X"00",X"25",X"9D",X"00",X"26",X"9D",X"00",
		X"27",X"9D",X"00",X"28",X"9D",X"00",X"29",X"9D",X"00",X"2A",X"9D",X"00",X"2B",X"9D",X"00",X"2C",
		X"9D",X"00",X"2D",X"9D",X"00",X"2E",X"9D",X"00",X"2F",X"8D",X"00",X"14",X"E8",X"D0",X"C1",X"8D",
		X"00",X"16",X"AD",X"00",X"08",X"29",X"10",X"D0",X"08",X"A9",X"20",X"8D",X"40",X"18",X"4C",X"CB",
		X"7B",X"A9",X"01",X"8D",X"00",X"20",X"A9",X"E4",X"8D",X"01",X"20",X"A9",X"20",X"8D",X"02",X"20",
		X"8D",X"03",X"20",X"8D",X"02",X"28",X"8D",X"03",X"28",X"A9",X"01",X"85",X"C4",X"85",X"CD",X"A9",
		X"FE",X"8D",X"24",X"18",X"E8",X"8D",X"26",X"18",X"A2",X"1D",X"A0",X"00",X"BD",X"7D",X"7B",X"9D",
		X"1C",X"03",X"A9",X"05",X"9D",X"FE",X"02",X"BD",X"7E",X"7B",X"9D",X"1D",X"03",X"BD",X"7F",X"7B",
		X"9D",X"1E",X"03",X"C8",X"CA",X"CA",X"CA",X"10",X"E3",X"20",X"1F",X"53",X"4C",X"00",X"50",X"1E",
		X"1C",X"38",X"2E",X"34",X"24",X"28",X"1E",X"1C",X"1C",X"1E",X"3A",X"3C",X"2A",X"1E",X"40",X"2A",
		X"18",X"1E",X"2C",X"00",X"24",X"16",X"1C",X"32",X"38",X"38",X"22",X"28",X"38",X"E3",X"A0",X"02",
		X"38",X"08",X"88",X"84",X"09",X"18",X"65",X"09",X"28",X"AA",X"08",X"86",X"08",X"B5",X"00",X"4A",
		X"4A",X"4A",X"4A",X"28",X"20",X"29",X"7A",X"A5",X"09",X"D0",X"01",X"18",X"A6",X"08",X"B5",X"00",
		X"20",X"29",X"7A",X"A6",X"08",X"CA",X"C6",X"09",X"10",X"E0",X"60",X"A2",X"11",X"9A",X"8A",X"85",
		X"00",X"A0",X"00",X"A2",X"01",X"C8",X"B9",X"00",X"00",X"D0",X"21",X"E8",X"D0",X"F7",X"BA",X"8A",
		X"8D",X"00",X"14",X"C8",X"59",X"00",X"00",X"D0",X"13",X"8A",X"A2",X"00",X"96",X"00",X"C8",X"D0",
		X"05",X"0A",X"A2",X"00",X"B0",X"4E",X"AA",X"9A",X"96",X"00",X"D0",X"D7",X"AA",X"8A",X"A0",X"82",
		X"29",X"0F",X"F0",X"02",X"A0",X"12",X"8A",X"A2",X"82",X"29",X"F0",X"F0",X"02",X"A2",X"12",X"98",
		X"9A",X"AA",X"8E",X"20",X"18",X"A2",X"A8",X"8E",X"21",X"18",X"A0",X"0C",X"A2",X"64",X"2C",X"00",
		X"08",X"30",X"FB",X"2C",X"00",X"08",X"10",X"FB",X"8D",X"00",X"14",X"CA",X"D0",X"F0",X"C0",X"05",
		X"D0",X"03",X"8E",X"21",X"18",X"88",X"D0",X"E4",X"4A",X"B0",X"03",X"BA",X"D0",X"D4",X"8D",X"00",
		X"14",X"4C",X"3E",X"7C",X"A2",X"7F",X"9A",X"A2",X"00",X"8A",X"95",X"00",X"E8",X"D0",X"FB",X"A8",
		X"A9",X"01",X"85",X"01",X"A2",X"11",X"B1",X"00",X"D0",X"27",X"8A",X"91",X"00",X"51",X"00",X"D0",
		X"20",X"8A",X"0A",X"AA",X"90",X"F4",X"C8",X"D0",X"EB",X"8D",X"00",X"14",X"E6",X"01",X"A6",X"01",
		X"E0",X"04",X"90",X"E0",X"A9",X"20",X"E0",X"20",X"90",X"D8",X"E0",X"30",X"90",X"D6",X"4C",X"01",
		X"7D",X"A6",X"01",X"E0",X"20",X"85",X"02",X"90",X"03",X"8A",X"E9",X"1C",X"4A",X"4A",X"29",X"07",
		X"A8",X"A5",X"02",X"84",X"00",X"85",X"01",X"A9",X"01",X"85",X"02",X"A2",X"A8",X"A0",X"82",X"A5",
		X"00",X"D0",X"08",X"A5",X"01",X"29",X"0F",X"F0",X"02",X"A0",X"12",X"8E",X"21",X"18",X"8C",X"20",
		X"18",X"A9",X"09",X"C0",X"12",X"F0",X"02",X"A9",X"01",X"A8",X"A2",X"00",X"2C",X"00",X"08",X"30",
		X"FB",X"2C",X"00",X"08",X"10",X"FB",X"8D",X"00",X"14",X"CA",X"D0",X"F0",X"88",X"D0",X"ED",X"8E",
		X"21",X"18",X"A0",X"09",X"2C",X"00",X"08",X"30",X"FB",X"2C",X"00",X"08",X"10",X"FB",X"8D",X"00",
		X"14",X"CA",X"D0",X"F0",X"88",X"D0",X"ED",X"A5",X"00",X"D0",X"08",X"A5",X"01",X"4A",X"4A",X"4A",
		X"4A",X"85",X"01",X"C6",X"02",X"F0",X"A4",X"C6",X"00",X"10",X"9C",X"8D",X"00",X"14",X"4C",X"FB",
		X"7C",X"A9",X"00",X"A8",X"AA",X"85",X"08",X"A9",X"30",X"85",X"09",X"A9",X"08",X"85",X"0A",X"A9",
		X"FF",X"51",X"08",X"C8",X"D0",X"FB",X"E6",X"09",X"8D",X"00",X"14",X"C6",X"0A",X"D0",X"F2",X"95",
		X"3D",X"E8",X"A5",X"09",X"C9",X"40",X"D0",X"04",X"A9",X"50",X"85",X"09",X"C9",X"80",X"90",X"D9",
		X"A2",X"FF",X"AD",X"00",X"08",X"29",X"20",X"D0",X"01",X"E8",X"86",X"0C",X"A2",X"00",X"18",X"BD",
		X"87",X"7D",X"30",X"40",X"29",X"1F",X"A8",X"BD",X"88",X"7D",X"99",X"60",X"18",X"A0",X"08",X"2C",
		X"00",X"18",X"10",X"07",X"88",X"10",X"F8",X"A9",X"54",X"D0",X"28",X"BD",X"87",X"7D",X"0A",X"A8",
		X"10",X"0D",X"AD",X"10",X"18",X"DD",X"89",X"7D",X"F0",X"04",X"A9",X"4C",X"D0",X"15",X"E8",X"98",
		X"0A",X"10",X"09",X"AD",X"18",X"18",X"DD",X"89",X"7D",X"D0",X"06",X"E8",X"E8",X"E8",X"4C",X"3E",
		X"7D",X"A9",X"48",X"38",X"4C",X"F4",X"7D",X"40",X"00",X"00",X"61",X"7F",X"00",X"7F",X"42",X"00",
		X"00",X"63",X"00",X"00",X"00",X"44",X"00",X"00",X"65",X"00",X"00",X"00",X"46",X"00",X"00",X"67",
		X"00",X"00",X"00",X"48",X"00",X"00",X"69",X"01",X"00",X"01",X"4A",X"80",X"80",X"6B",X"00",X"7F",
		X"00",X"6C",X"10",X"10",X"00",X"72",X"00",X"3F",X"00",X"78",X"00",X"00",X"80",X"79",X"00",X"3F",
		X"00",X"77",X"00",X"7F",X"00",X"73",X"00",X"00",X"80",X"40",X"00",X"00",X"61",X"5A",X"00",X"5A",
		X"42",X"00",X"00",X"63",X"A6",X"00",X"A6",X"44",X"FF",X"FF",X"65",X"7F",X"FF",X"7F",X"46",X"FF",
		X"FF",X"67",X"7F",X"FF",X"7F",X"48",X"00",X"00",X"69",X"01",X"00",X"01",X"4A",X"00",X"00",X"6B",
		X"01",X"B4",X"A6",X"FF",X"B0",X"02",X"A9",X"00",X"85",X"0D",X"A5",X"3D",X"F0",X"0A",X"A9",X"F0",
		X"A2",X"A2",X"8D",X"20",X"18",X"8E",X"21",X"18",X"A9",X"02",X"85",X"00",X"A9",X"00",X"85",X"01",
		X"A2",X"28",X"2C",X"00",X"08",X"10",X"FB",X"2C",X"00",X"08",X"30",X"FB",X"CA",X"10",X"F3",X"2C",
		X"00",X"08",X"50",X"FB",X"8D",X"00",X"14",X"A9",X"00",X"85",X"02",X"A9",X"20",X"85",X"03",X"24",
		X"0C",X"30",X"36",X"20",X"6A",X"7A",X"A9",X"81",X"AA",X"A0",X"00",X"20",X"8E",X"7A",X"A9",X"00",
		X"20",X"63",X"7A",X"20",X"6A",X"7A",X"A9",X"7F",X"AA",X"A0",X"00",X"20",X"8E",X"7A",X"A9",X"02",
		X"20",X"63",X"7A",X"A6",X"0C",X"BC",X"CA",X"7F",X"A9",X"20",X"91",X"02",X"88",X"88",X"B9",X"CE",
		X"7F",X"91",X"02",X"88",X"10",X"F8",X"4C",X"2A",X"7F",X"A9",X"37",X"A2",X"0A",X"20",X"5A",X"7A",
		X"20",X"6A",X"7A",X"A9",X"82",X"A2",X"A7",X"20",X"90",X"7A",X"A9",X"33",X"A2",X"F0",X"20",X"5A",
		X"7A",X"20",X"6A",X"7A",X"A9",X"D3",X"A2",X"13",X"20",X"90",X"7A",X"A2",X"0F",X"AD",X"00",X"0A",
		X"49",X"FF",X"85",X"0B",X"AD",X"00",X"0C",X"49",X"FF",X"48",X"86",X"0A",X"29",X"01",X"20",X"2F",
		X"7A",X"A6",X"0A",X"46",X"0B",X"68",X"6A",X"CA",X"10",X"EF",X"20",X"6A",X"7A",X"A9",X"FB",X"A2",
		X"1D",X"20",X"90",X"7A",X"A9",X"01",X"20",X"2F",X"7A",X"AD",X"00",X"0C",X"29",X"10",X"4A",X"4A",
		X"4A",X"4A",X"69",X"01",X"20",X"2F",X"7A",X"AD",X"00",X"0C",X"29",X"0C",X"4A",X"4A",X"AA",X"BD",
		X"C6",X"7F",X"20",X"2F",X"7A",X"A2",X"16",X"86",X"0B",X"A2",X"07",X"B5",X"3D",X"F0",X"29",X"85",
		X"00",X"86",X"0A",X"20",X"6A",X"7A",X"A6",X"0B",X"8A",X"38",X"E9",X"08",X"85",X"0B",X"A9",X"A0",
		X"20",X"90",X"7A",X"A5",X"0A",X"20",X"2F",X"7A",X"A9",X"06",X"A2",X"00",X"20",X"90",X"7A",X"A9",
		X"00",X"A0",X"01",X"20",X"A0",X"7B",X"A6",X"0A",X"CA",X"10",X"D0",X"20",X"6A",X"7A",X"A9",X"60",
		X"A2",X"16",X"20",X"90",X"7A",X"A5",X"0D",X"F0",X"0E",X"38",X"E9",X"36",X"0A",X"A8",X"B9",X"F0",
		X"33",X"BE",X"F1",X"33",X"20",X"6E",X"7A",X"20",X"1D",X"7A",X"8D",X"00",X"12",X"24",X"0C",X"10",
		X"4D",X"20",X"B9",X"7F",X"D0",X"4D",X"8D",X"2B",X"18",X"A0",X"00",X"AD",X"28",X"18",X"29",X"7F",
		X"4A",X"90",X"01",X"C8",X"09",X"00",X"D0",X"F8",X"AD",X"00",X"08",X"29",X"0F",X"49",X"0F",X"4A",
		X"90",X"01",X"C8",X"09",X"00",X"D0",X"F8",X"C4",X"10",X"F0",X"08",X"A9",X"A7",X"90",X"08",X"A2",
		X"80",X"D0",X"06",X"A9",X"00",X"F0",X"02",X"A2",X"20",X"84",X"10",X"8D",X"23",X"18",X"8E",X"22",
		X"18",X"AD",X"00",X"08",X"29",X"10",X"D0",X"03",X"4C",X"3C",X"7D",X"4C",X"CC",X"7A",X"20",X"B9",
		X"7F",X"F0",X"F5",X"E6",X"0C",X"A5",X"0C",X"29",X"FC",X"F0",X"ED",X"A9",X"00",X"8D",X"00",X"14",
		X"8D",X"40",X"18",X"8D",X"60",X"18",X"8D",X"20",X"18",X"AD",X"00",X"18",X"AD",X"18",X"18",X"AD",
		X"10",X"18",X"A9",X"01",X"8D",X"40",X"18",X"A2",X"1F",X"18",X"9D",X"60",X"18",X"2A",X"CA",X"10",
		X"F9",X"20",X"B9",X"7F",X"F0",X"D5",X"4C",X"CC",X"7A",X"AD",X"00",X"08",X"A8",X"45",X"13",X"25",
		X"13",X"84",X"13",X"29",X"20",X"60",X"01",X"04",X"05",X"06",X"0D",X"11",X"17",X"2D",X"40",X"80",
		X"80",X"1E",X"00",X"1E",X"FF",X"02",X"FF",X"E3",X"40",X"80",X"0F",X"51",X"F1",X"4F",X"12",X"E0",
		X"00",X"20",X"F1",X"4F",X"16",X"A0",X"E0",X"51",X"00",X"20",X"18",X"A0",X"00",X"C0",X"1A",X"A0",
		X"00",X"C0",X"1C",X"A0",X"00",X"C0",X"EF",X"40",X"00",X"C0",X"8F",X"55",X"CC",X"7A",X"CC",X"7A");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
