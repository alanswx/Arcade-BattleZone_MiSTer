

`define OP_VCTR    3'b000
`define OP_HALT    3'b001
`define OP_SVEC    3'b010
`define OP_STORE   3'b011
`define OP_CNTR    3'b100
`define OP_JSR     3'b101
`define OP_RTS     3'b110
`define OP_JMP     3'b111
