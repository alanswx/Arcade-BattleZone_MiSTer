
`define BRAM_PROG_RAM 3'b000
`define BRAM_VECTOR   3'b001
`define BRAM_PROG_ROM 3'b010
`define BRAM_POKEY 3'b011
`define BRAM_MATH 3'b100
