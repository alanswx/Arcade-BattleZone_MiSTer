module auxPCB
  (

   );

endmodule: auxPCB
