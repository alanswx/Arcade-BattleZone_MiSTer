library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity C:\Users\hp\Desktop\F15_18545_BattleZone-master\rtl\roms\vec is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of C:\Users\hp\Desktop\F15_18545_BattleZone-master\rtl\roms\vec is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"7A",X"00",X"C0",X"0B",X"A8",X"65",X"A8",X"82",X"A8",X"C1",X"A8",X"E2",X"A8",
		X"F9",X"A8",X"17",X"A9",X"34",X"A9",X"40",X"00",X"00",X"00",X"E0",X"1F",X"20",X"60",X"18",X"5C",
		X"28",X"00",X"50",X"60",X"00",X"00",X"20",X"60",X"E0",X"1F",X"20",X"60",X"20",X"00",X"C0",X"7F",
		X"C0",X"1F",X"00",X"00",X"40",X"00",X"80",X"60",X"C0",X"1F",X"40",X"60",X"00",X"00",X"20",X"00",
		X"20",X"00",X"C0",X"7F",X"20",X"00",X"E0",X"1F",X"E0",X"1F",X"40",X"60",X"F0",X"1F",X"40",X"60",
		X"F0",X"1F",X"60",X"60",X"A0",X"00",X"30",X"00",X"F4",X"1F",X"05",X"E0",X"E0",X"5A",X"FC",X"5A",
		X"FA",X"5A",X"FD",X"1F",X"F4",X"FF",X"03",X"00",X"F4",X"FF",X"F7",X"1F",X"0C",X"E0",X"FD",X"1F",
		X"0C",X"E0",X"03",X"00",X"0C",X"E0",X"09",X"00",X"0C",X"E0",X"E3",X"46",X"E0",X"46",X"FE",X"46",
		X"0C",X"00",X"F5",X"FF",X"03",X"00",X"F3",X"5F",X"FC",X"1F",X"F1",X"5F",X"5B",X"5C",X"F5",X"1F",
		X"FB",X"5F",X"F3",X"1F",X"FE",X"5F",X"F1",X"1F",X"06",X"40",X"03",X"00",X"1B",X"00",X"A0",X"5E",
		X"FF",X"1F",X"06",X"A0",X"0B",X"00",X"06",X"A0",X"FF",X"1F",X"FC",X"BF",X"02",X"00",X"FF",X"BF",
		X"09",X"4A",X"FD",X"1F",X"FD",X"BF",X"03",X"00",X"01",X"A0",X"01",X"00",X"FD",X"BF",X"A0",X"43",
		X"01",X"00",X"01",X"40",X"6A",X"1F",X"07",X"00",X"00",X"C0",X"00",X"00",X"20",X"00",X"30",X"00",
		X"40",X"60",X"D0",X"1F",X"20",X"60",X"30",X"00",X"E0",X"1F",X"F0",X"1F",X"20",X"60",X"20",X"00",
		X"40",X"60",X"C0",X"1F",X"A0",X"60",X"20",X"00",X"80",X"7F",X"20",X"00",X"E0",X"7F",X"E0",X"1F",
		X"C0",X"1F",X"E0",X"1F",X"60",X"60",X"00",X"00",X"80",X"00",X"20",X"00",X"A0",X"60",X"E0",X"1F",
		X"00",X"00",X"00",X"C0",X"20",X"00",X"00",X"00",X"00",X"00",X"40",X"60",X"E0",X"1F",X"00",X"00",
		X"20",X"00",X"C0",X"7F",X"00",X"00",X"40",X"00",X"20",X"00",X"40",X"60",X"E0",X"1F",X"C0",X"1F",
		X"E0",X"1F",X"60",X"60",X"20",X"00",X"20",X"60",X"20",X"00",X"C0",X"7F",X"00",X"00",X"20",X"60",
		X"E0",X"1F",X"20",X"60",X"10",X"00",X"20",X"60",X"F0",X"1F",X"20",X"60",X"E0",X"1F",X"A0",X"7F",
		X"20",X"00",X"60",X"00",X"20",X"00",X"40",X"60",X"E0",X"1F",X"40",X"60",X"10",X"00",X"A0",X"1F",
		X"F0",X"1F",X"20",X"60",X"10",X"00",X"20",X"60",X"D0",X"1F",X"00",X"00",X"08",X"00",X"60",X"60",
		X"18",X"00",X"C0",X"7F",X"10",X"00",X"20",X"60",X"F0",X"1F",X"40",X"60",X"E8",X"1F",X"E0",X"7F",
		X"28",X"00",X"E0",X"7F",X"F0",X"1F",X"40",X"00",X"00",X"00",X"20",X"60",X"E0",X"1F",X"00",X"00",
		X"00",X"C0",X"20",X"00",X"00",X"00",X"E0",X"1F",X"40",X"60",X"20",X"00",X"C0",X"1F",X"E0",X"1F",
		X"80",X"60",X"00",X"00",X"A0",X"00",X"20",X"00",X"60",X"60",X"E0",X"1F",X"20",X"60",X"20",X"00",
		X"E0",X"1F",X"20",X"00",X"20",X"60",X"C0",X"1F",X"20",X"60",X"00",X"00",X"20",X"00",X"40",X"00",
		X"C0",X"7F",X"E0",X"1F",X"20",X"00",X"20",X"00",X"20",X"60",X"E0",X"1F",X"20",X"60",X"E0",X"1F",
		X"00",X"00",X"00",X"C0",X"20",X"00",X"00",X"00",X"20",X"00",X"40",X"60",X"C0",X"1F",X"20",X"60",
		X"00",X"00",X"20",X"00",X"40",X"00",X"C0",X"7F",X"E0",X"1F",X"20",X"00",X"10",X"00",X"20",X"60",
		X"D0",X"1F",X"60",X"60",X"00",X"00",X"80",X"00",X"20",X"00",X"A0",X"60",X"E0",X"1F",X"00",X"00",
		X"00",X"C0",X"20",X"00",X"00",X"00",X"00",X"00",X"40",X"60",X"E0",X"1F",X"E0",X"60",X"30",X"00",
		X"E0",X"7F",X"E0",X"1F",X"C0",X"7F",X"F0",X"1F",X"60",X"00",X"40",X"00",X"60",X"60",X"D8",X"1F",
		X"40",X"60",X"18",X"54",X"60",X"00",X"40",X"60",X"F9",X"1F",X"03",X"60",X"05",X"00",X"05",X"60",
		X"FA",X"1F",X"03",X"60",X"08",X"00",X"05",X"60",X"A0",X"1F",X"00",X"00",X"00",X"C0",X"60",X"00",
		X"00",X"00",X"A0",X"1F",X"40",X"60",X"40",X"00",X"60",X"60",X"C0",X"1F",X"40",X"60",X"00",X"00",
		X"40",X"00",X"40",X"00",X"80",X"7F",X"E0",X"1F",X"40",X"00",X"20",X"00",X"40",X"60",X"C0",X"1F",
		X"80",X"60",X"20",X"00",X"C0",X"1F",X"10",X"00",X"40",X"60",X"D0",X"1F",X"20",X"60",X"30",X"00",
		X"E0",X"1F",X"D0",X"1F",X"60",X"60",X"00",X"C0",X"00",X"00",X"C0",X"00",X"20",X"00",X"E0",X"60",
		X"E0",X"1F",X"40",X"60",X"10",X"00",X"E0",X"1F",X"30",X"00",X"40",X"60",X"C0",X"1F",X"00",X"00",
		X"00",X"C0",X"C0",X"48",X"C4",X"44",X"C4",X"5C",X"C0",X"58",X"18",X"44",X"C8",X"40",X"04",X"5C",
		X"00",X"C0",X"C0",X"4C",X"C6",X"40",X"C2",X"5E",X"C0",X"5E",X"DE",X"5E",X"DA",X"40",X"06",X"40",
		X"C2",X"5E",X"C0",X"5E",X"DE",X"5E",X"DA",X"40",X"93",X"E9",X"C0",X"4C",X"C8",X"40",X"18",X"54",
		X"D6",X"E9",X"C0",X"4C",X"C4",X"40",X"C4",X"5C",X"C0",X"5C",X"DC",X"5C",X"DC",X"40",X"93",X"E9",
		X"C8",X"40",X"18",X"40",X"C0",X"4C",X"C8",X"40",X"1E",X"5A",X"DA",X"40",X"0C",X"5A",X"00",X"C0",
		X"C0",X"4C",X"C8",X"40",X"C0",X"5C",X"1C",X"5C",X"C4",X"40",X"C0",X"5C",X"92",X"E9",X"C0",X"4C",
		X"00",X"5A",X"C8",X"40",X"00",X"46",X"EF",X"E9",X"C8",X"40",X"18",X"4C",X"C8",X"40",X"1C",X"40",
		X"C0",X"54",X"08",X"40",X"00",X"C0",X"00",X"44",X"C4",X"5C",X"C4",X"40",X"B4",X"E9",X"C0",X"4C",
		X"06",X"40",X"DA",X"5A",X"C6",X"5A",X"06",X"40",X"00",X"C0",X"00",X"4C",X"C0",X"54",X"D6",X"E9",
		X"C0",X"4C",X"C4",X"5C",X"C4",X"44",X"EF",X"E9",X"C0",X"4C",X"C8",X"54",X"B4",X"E9",X"C0",X"4C",
		X"C8",X"40",X"C0",X"54",X"D8",X"40",X"0C",X"40",X"00",X"C0",X"C0",X"4C",X"C8",X"40",X"C0",X"5A",
		X"D8",X"40",X"66",X"E9",X"C0",X"4C",X"C8",X"40",X"C0",X"58",X"DC",X"5C",X"DC",X"40",X"04",X"44",
		X"C4",X"5C",X"D7",X"E9",X"C0",X"4C",X"C8",X"40",X"C0",X"5A",X"D8",X"40",X"02",X"40",X"C6",X"5A",
		X"D7",X"E9",X"C8",X"40",X"C0",X"46",X"D8",X"40",X"C0",X"46",X"C8",X"40",X"B5",X"E9",X"00",X"4C",
		X"76",X"E9",X"00",X"4C",X"C0",X"54",X"C8",X"40",X"C0",X"4C",X"04",X"54",X"00",X"C0",X"00",X"4C",
		X"C4",X"54",X"C4",X"4C",X"B5",X"E9",X"00",X"4C",X"C0",X"54",X"C4",X"44",X"C4",X"5C",X"B4",X"E9",
		X"C8",X"4C",X"18",X"40",X"C8",X"54",X"F0",X"E9",X"04",X"40",X"C0",X"48",X"DC",X"44",X"08",X"40",
		X"DC",X"5C",X"08",X"58",X"00",X"C0",X"00",X"4C",X"C8",X"40",X"D8",X"54",X"D6",X"E9",X"04",X"4C",
		X"78",X"E9",X"00",X"4C",X"C8",X"40",X"C0",X"5A",X"D8",X"40",X"C0",X"5A",X"C8",X"40",X"04",X"40",
		X"00",X"C0",X"00",X"4C",X"C8",X"40",X"C0",X"54",X"D8",X"40",X"00",X"46",X"C8",X"40",X"04",X"5A",
		X"00",X"C0",X"00",X"4C",X"C0",X"5A",X"C8",X"40",X"00",X"46",X"EF",X"E9",X"00",X"46",X"C8",X"40",
		X"C0",X"5A",X"D8",X"40",X"C0",X"4C",X"0C",X"54",X"00",X"C0",X"00",X"4C",X"C8",X"40",X"C0",X"54",
		X"04",X"40",X"00",X"C0",X"C0",X"4C",X"DA",X"E9",X"08",X"46",X"D8",X"40",X"C0",X"46",X"EE",X"E9",
		X"93",X"A9",X"8F",X"A9",X"CF",X"A9",X"D1",X"A9",X"D9",X"A9",X"E1",X"A9",X"A9",X"A9",X"E6",X"A9",
		X"ED",X"A9",X"F2",X"A9",X"F4",X"A9",X"41",X"A9",X"49",X"A9",X"55",X"A9",X"59",X"A9",X"60",X"A9",
		X"62",X"A9",X"68",X"A9",X"6F",X"A9",X"74",X"A9",X"7B",X"A9",X"7F",X"A9",X"85",X"A9",X"88",X"A9",
		X"8C",X"A9",X"8F",X"A9",X"95",X"A9",X"9A",X"A9",X"A2",X"A9",X"A9",X"A9",X"AF",X"A9",X"B1",X"A9",
		X"B7",X"A9",X"BB",X"A9",X"C0",X"A9",X"C4",X"A9",X"CB",X"A9",X"93",X"A9",X"D6",X"A9",X"2A",X"AA",
		X"33",X"AA",X"00",X"C0",X"00",X"42",X"C0",X"48",X"C4",X"42",X"C4",X"5E",X"C0",X"58",X"DC",X"5E",
		X"DC",X"42",X"00",X"C0",X"22",X"AA",X"01",X"00",X"0B",X"00",X"DD",X"40",X"C0",X"47",X"C3",X"40",
		X"ED",X"1F",X"0D",X"00",X"00",X"C0",X"22",X"AA",X"01",X"00",X"05",X"00",X"C0",X"47",X"C3",X"40",
		X"C0",X"5D",X"DD",X"40",X"F3",X"1F",X"13",X"00",X"00",X"C0",X"00",X"00",X"C0",X"1F",X"00",X"00",
		X"00",X"E0",X"C0",X"1F",X"C0",X"1F",X"00",X"00",X"00",X"E0",X"C0",X"1F",X"40",X"00",X"00",X"00",
		X"00",X"E0",X"20",X"00",X"60",X"00",X"00",X"00",X"00",X"E0",X"E0",X"1F",X"40",X"00",X"00",X"00",
		X"00",X"E0",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"60",X"00",X"20",X"00",X"00",X"00",
		X"00",X"E0",X"60",X"00",X"E0",X"1F",X"00",X"00",X"00",X"E0",X"E0",X"1F",X"80",X"1F",X"00",X"00",
		X"00",X"E0",X"20",X"00",X"A0",X"1F",X"00",X"00",X"00",X"E0",X"00",X"C0",X"40",X"80",X"51",X"1F",
		X"00",X"00",X"64",X"00",X"00",X"60",X"19",X"00",X"B5",X"1F",X"E7",X"1F",X"00",X"60",X"00",X"00",
		X"96",X"60",X"19",X"00",X"00",X"60",X"64",X"00",X"00",X"00",X"19",X"00",X"00",X"60",X"00",X"00",
		X"6A",X"7F",X"E7",X"1F",X"00",X"60",X"19",X"00",X"4B",X"00",X"64",X"00",X"00",X"60",X"00",X"C0",
		X"40",X"80",X"51",X"1F",X"00",X"00",X"64",X"00",X"00",X"E0",X"28",X"00",X"00",X"60",X"00",X"00",
		X"DD",X"1F",X"D8",X"1F",X"D8",X"FF",X"00",X"00",X"96",X"E0",X"28",X"00",X"D8",X"FF",X"46",X"00",
		X"00",X"00",X"28",X"00",X"28",X"E0",X"00",X"00",X"6A",X"FF",X"D8",X"1F",X"28",X"E0",X"00",X"00",
		X"23",X"00",X"28",X"00",X"00",X"60",X"64",X"00",X"00",X"E0",X"00",X"C0",X"40",X"80",X"3C",X"01",
		X"44",X"00",X"FC",X"40",X"C4",X"1F",X"C4",X"1F",X"E0",X"5C",X"44",X"00",X"C4",X"1F",X"FC",X"40",
		X"00",X"00",X"44",X"00",X"34",X"00",X"DC",X"BF",X"08",X"00",X"24",X"00",X"E0",X"44",X"F0",X"1F",
		X"24",X"00",X"CC",X"1F",X"DC",X"BF",X"00",X"C0",X"DD",X"43",X"03",X"00",X"09",X"C0",X"06",X"00",
		X"03",X"C0",X"F7",X"1F",X"24",X"C0",X"DD",X"5D",X"00",X"00",X"DC",X"DF",X"09",X"46",X"00",X"00",
		X"15",X"C0",X"FD",X"1F",X"00",X"C0",X"00",X"00",X"F7",X"DF",X"F7",X"1F",X"1B",X"00",X"00",X"C0",
		X"B4",X"AA",X"40",X"80",X"32",X"00",X"9C",X"1F",X"00",X"00",X"B5",X"DF",X"9C",X"1F",X"23",X"00",
		X"64",X"00",X"28",X"C0",X"64",X"00",X"9C",X"DF",X"19",X"00",X"FA",X"00",X"83",X"1F",X"6A",X"DF",
		X"CE",X"1F",X"64",X"C0",X"00",X"C0",X"00",X"00",X"50",X"C0",X"CE",X"1F",X"24",X"1F",X"CE",X"1F",
		X"41",X"C0",X"96",X"00",X"9C",X"1F",X"D3",X"1F",X"00",X"C0",X"91",X"00",X"E7",X"1F",X"2D",X"00",
		X"6A",X"DF",X"1E",X"00",X"E1",X"00",X"B5",X"1F",X"B5",X"DF",X"19",X"00",X"FA",X"00",X"5F",X"00",
		X"0A",X"C0",X"A1",X"1F",X"F6",X"1F",X"3C",X"00",X"64",X"C0",X"00",X"C0",X"3C",X"00",X"64",X"C0",
		X"2D",X"00",X"9C",X"1F",X"97",X"1F",X"00",X"C0",X"F6",X"1F",X"ED",X"1E",X"5F",X"00",X"97",X"DF",
		X"83",X"1F",X"88",X"1F",X"0A",X"00",X"CE",X"DF",X"F6",X"1F",X"32",X"00",X"88",X"1F",X"7E",X"DF",
		X"BA",X"1F",X"31",X"01",X"FB",X"1F",X"A6",X"DF",X"9C",X"1F",X"BE",X"00",X"74",X"1F",X"2D",X"C0",
		X"F0",X"00",X"6E",X"00",X"D8",X"1F",X"00",X"C0",X"00",X"C0",X"00",X"00",X"69",X"C0",X"38",X"1F",
		X"29",X"1F",X"6A",X"1F",X"B0",X"DF",X"86",X"01",X"65",X"1F",X"CE",X"1F",X"00",X"C0",X"32",X"00",
		X"00",X"00",X"19",X"00",X"AB",X"DF",X"27",X"01",X"78",X"00",X"73",X"00",X"88",X"DF",X"0F",X"00",
		X"AF",X"00",X"7E",X"1F",X"C9",X"DF",X"E7",X"1F",X"E0",X"01",X"00",X"00",X"46",X"C0",X"69",X"00",
		X"3D",X"1F",X"C4",X"1F",X"19",X"C0",X"55",X"00",X"4B",X"C0",X"00",X"C0",X"41",X"00",X"F1",X"DF",
		X"D8",X"1F",X"32",X"00",X"E7",X"1F",X"DD",X"DF",X"2F",X"1E",X"D8",X"1F",X"64",X"00",X"69",X"C0",
		X"60",X"1F",X"B0",X"1F",X"3C",X"00",X"E7",X"DF",X"C4",X"1F",X"F6",X"DF",X"A2",X"1E",X"06",X"1F",
		X"3C",X"00",X"DD",X"DF",X"C4",X"1F",X"D8",X"DF",X"90",X"01",X"8D",X"1F",X"E2",X"1F",X"DD",X"DF",
		X"00",X"C0",X"BA",X"1F",X"32",X"C0",X"1E",X"00",X"9C",X"1F",X"28",X"00",X"32",X"C0",X"EC",X"1F",
		X"DB",X"01",X"CE",X"1F",X"CE",X"DF",X"58",X"02",X"87",X"00",X"CE",X"1F",X"0F",X"C0",X"AC",X"1E",
		X"0F",X"00",X"92",X"1F",X"5F",X"C0",X"00",X"C0",X"4B",X"00",X"73",X"C0",X"8D",X"1F",X"A6",X"1F",
		X"28",X"00",X"E7",X"DF",X"BA",X"1F",X"21",X"1D",X"F1",X"1F",X"BF",X"DF",X"00",X"C0",X"2D",X"00",
		X"AB",X"DF",X"A1",X"1F",X"32",X"00",X"32",X"00",X"23",X"C0",X"F1",X"1F",X"57",X"03",X"3C",X"00",
		X"E2",X"DF",X"1E",X"00",X"50",X"C0",X"00",X"C0",X"C9",X"AA",X"DB",X"AA",X"F6",X"AA",X"15",X"AB",
		X"36",X"AB",X"51",X"AB",X"64",X"AB",X"6F",X"AB",X"00",X"C0",X"40",X"80",X"00",X"71",X"08",X"02",
		X"08",X"02",X"10",X"62",X"40",X"80",X"F8",X"1D",X"F8",X"1D",X"20",X"60",X"88",X"00",X"08",X"00",
		X"00",X"00",X"FF",X"E3",X"FF",X"02",X"00",X"E0",X"00",X"00",X"01",X"FC",X"01",X"1D",X"00",X"E0",
		X"FF",X"02",X"FF",X"E2",X"00",X"1F",X"00",X"E1",X"01",X"1E",X"01",X"FE",X"00",X"02",X"00",X"FE",
		X"FF",X"00",X"00",X"E1",X"01",X"1D",X"FF",X"E2",X"FF",X"02",X"00",X"00",X"01",X"1D",X"01",X"FD",
		X"FF",X"00",X"00",X"FF",X"00",X"02",X"00",X"E2",X"01",X"1E",X"FF",X"E1",X"00",X"1F",X"00",X"FF",
		X"FF",X"02",X"01",X"FD",X"40",X"80",X"18",X"5C",X"EF",X"40",X"1F",X"42",X"D3",X"40",X"01",X"42",
		X"AB",X"40",X"1F",X"42",X"97",X"40",X"01",X"42",X"67",X"40",X"1F",X"42",X"5B",X"40",X"01",X"42",
		X"23",X"40",X"00",X"C0",X"92",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"01",X"01",X"01",X"02",
		X"02",X"02",X"02",X"02",X"02",X"03",X"03",X"03",X"03",X"03",X"03",X"03",X"04",X"04",X"04",X"04",
		X"04",X"04",X"05",X"05",X"05",X"05",X"05",X"05",X"06",X"06",X"06",X"06",X"06",X"06",X"06",X"07",
		X"07",X"07",X"07",X"07",X"07",X"08",X"08",X"08",X"08",X"08",X"08",X"08",X"09",X"09",X"09",X"09",
		X"09",X"09",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0E",X"0E",
		X"0E",X"0E",X"0E",X"0E",X"0E",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"10",X"10",X"10",X"10",
		X"10",X"10",X"10",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"12",X"12",X"12",X"12",X"12",
		X"12",X"12",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"13",X"14",X"14",X"14",X"14",X"14",X"14",
		X"14",X"14",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"15",X"16",X"16",X"16",X"16",X"16",
		X"16",X"16",X"16",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"17",X"18",X"18",X"18",X"18",
		X"18",X"18",X"18",X"18",X"18",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"19",X"1A",
		X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1A",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",X"1B",
		X"1B",X"1B",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1D",X"1D",X"1D",
		X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1D",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",X"1E",
		X"1E",X"1E",X"1E",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"1F",X"20",
		X"20",X"20",X"20",X"20",X"20",X"D4",X"00",X"14",X"24",X"49",X"05",X"10",X"20",X"30",X"E6",X"38",
		X"05",X"39",X"55",X"39",X"36",X"39",X"55",X"3A",X"30",X"3A",X"0B",X"3A",X"E6",X"39",X"7A",X"3A",
		X"9F",X"3A",X"C4",X"3A",X"E9",X"3A",X"3B",X"3C",X"0E",X"3B",X"3F",X"3B",X"5A",X"3C",X"9B",X"3B",
		X"C0",X"3B",X"46",X"3B",X"0E",X"3B",X"C0",X"3B",X"9B",X"3B",X"8B",X"3C",X"D5",X"76",X"C0",X"3B",
		X"0A",X"3C",X"9B",X"3B",X"F1",X"3B",X"9B",X"3B",X"0A",X"3C",X"4E",X"77",X"CD",X"77",X"B0",X"3E",
		X"17",X"3F",X"00",X"00",X"00",X"00",X"28",X"3D",X"59",X"3D",X"8A",X"3D",X"BB",X"3D",X"EC",X"3D",
		X"1D",X"3E",X"4E",X"3E",X"7F",X"3E",X"1F",X"00",X"FE",X"00",X"FE",X"C0",X"FE",X"00",X"FE",X"00",
		X"02",X"C0",X"FE",X"00",X"02",X"00",X"02",X"C0",X"FE",X"00",X"02",X"00",X"FE",X"C0",X"FE",X"00",
		X"00",X"00",X"00",X"40",X"01",X"31",X"00",X"FE",X"00",X"FE",X"C0",X"FE",X"00",X"FE",X"00",X"02",
		X"C0",X"FE",X"00",X"02",X"00",X"02",X"C0",X"FE",X"00",X"02",X"00",X"FE",X"C0",X"FE",X"00",X"FE",
		X"00",X"FE",X"40",X"01",X"00",X"FE",X"00",X"02",X"40",X"01",X"00",X"02",X"00",X"02",X"40",X"01",
		X"00",X"02",X"00",X"FE",X"40",X"01",X"1F",X"D8",X"FF",X"D8",X"FF",X"D0",X"FF",X"D8",X"FF",X"D8",
		X"FF",X"F8",X"FF",X"D8",X"FF",X"28",X"00",X"F8",X"FF",X"D8",X"FF",X"28",X"00",X"D0",X"FF",X"50",
		X"00",X"00",X"00",X"E4",X"FF",X"91",X"20",X"FD",X"00",X"FE",X"C0",X"FE",X"20",X"FD",X"00",X"02",
		X"C0",X"FE",X"C8",X"03",X"00",X"02",X"C0",X"FE",X"C8",X"03",X"00",X"FE",X"C0",X"FE",X"00",X"FC",
		X"C8",X"FD",X"30",X"FF",X"00",X"FC",X"38",X"02",X"30",X"FF",X"E0",X"04",X"38",X"02",X"30",X"FF",
		X"E0",X"04",X"C8",X"FD",X"30",X"FF",X"58",X"FD",X"A8",X"FE",X"88",X"FF",X"58",X"FD",X"58",X"01",
		X"88",X"FF",X"A8",X"02",X"58",X"01",X"88",X"FF",X"A8",X"02",X"A8",X"FE",X"88",X"FF",X"00",X"FE",
		X"58",X"FF",X"30",X"00",X"00",X"FE",X"A8",X"00",X"30",X"00",X"80",X"FF",X"D8",X"FF",X"F8",X"FF",
		X"80",X"FF",X"28",X"00",X"F8",X"FF",X"80",X"00",X"28",X"00",X"D0",X"FF",X"80",X"00",X"D8",X"FF",
		X"D0",X"FF",X"60",X"04",X"28",X"00",X"F8",X"FF",X"60",X"04",X"28",X"00",X"D0",X"FF",X"60",X"04",
		X"D8",X"FF",X"F8",X"FF",X"60",X"04",X"D8",X"FF",X"D0",X"FF",X"00",X"FE",X"00",X"00",X"30",X"00",
		X"00",X"FE",X"00",X"00",X"50",X"00",X"25",X"00",X"FC",X"C8",X"FD",X"30",X"FF",X"00",X"FC",X"38",
		X"02",X"30",X"FF",X"68",X"FC",X"DC",X"FD",X"08",X"FF",X"68",X"FC",X"24",X"02",X"08",X"FF",X"D0",
		X"FC",X"EC",X"FD",X"E0",X"FE",X"D0",X"FC",X"14",X"02",X"E0",X"FE",X"25",X"18",X"FC",X"CC",X"FD",
		X"28",X"FF",X"18",X"FC",X"34",X"02",X"28",X"FF",X"80",X"FC",X"E0",X"FD",X"00",X"FF",X"80",X"FC",
		X"20",X"02",X"00",X"FF",X"E8",X"FC",X"F0",X"FD",X"D8",X"FE",X"E8",X"FC",X"10",X"02",X"D8",X"FE",
		X"25",X"34",X"FC",X"D4",X"FD",X"1C",X"FF",X"34",X"FC",X"2C",X"02",X"1C",X"FF",X"9C",X"FC",X"E4",
		X"FD",X"F4",X"FE",X"9C",X"FC",X"1C",X"02",X"F4",X"FE",X"04",X"FD",X"F8",X"FD",X"CC",X"FE",X"04",
		X"FD",X"08",X"02",X"CC",X"FE",X"25",X"4C",X"FC",X"D8",X"FD",X"14",X"FF",X"4C",X"FC",X"28",X"02",
		X"14",X"FF",X"B4",X"FC",X"E8",X"FD",X"EC",X"FE",X"B4",X"FC",X"18",X"02",X"EC",X"FE",X"20",X"FD",
		X"FC",X"FD",X"C4",X"FE",X"20",X"FD",X"04",X"02",X"C4",X"FE",X"25",X"E0",X"04",X"C8",X"FD",X"30",
		X"FF",X"E0",X"04",X"38",X"02",X"30",X"FF",X"80",X"04",X"DC",X"FD",X"08",X"FF",X"80",X"04",X"24",
		X"02",X"08",X"FF",X"20",X"04",X"EC",X"FD",X"E0",X"FE",X"20",X"04",X"14",X"02",X"E0",X"FE",X"25",
		X"C8",X"04",X"CC",X"FD",X"28",X"FF",X"C8",X"04",X"34",X"02",X"28",X"FF",X"68",X"04",X"E0",X"FD",
		X"00",X"FF",X"68",X"04",X"20",X"02",X"00",X"FF",X"08",X"04",X"F0",X"FD",X"D8",X"FE",X"08",X"04",
		X"10",X"02",X"D8",X"FE",X"25",X"B0",X"04",X"D4",X"FD",X"1C",X"FF",X"B0",X"04",X"2C",X"02",X"1C",
		X"FF",X"50",X"04",X"E4",X"FD",X"F4",X"FE",X"50",X"04",X"1C",X"02",X"F4",X"FE",X"F0",X"03",X"F8",
		X"FD",X"CC",X"FE",X"F0",X"03",X"08",X"02",X"CC",X"FE",X"25",X"98",X"04",X"D8",X"FD",X"14",X"FF",
		X"98",X"04",X"28",X"02",X"14",X"FF",X"38",X"04",X"E8",X"FD",X"EC",X"FE",X"38",X"04",X"18",X"02",
		X"EC",X"FE",X"D8",X"03",X"FC",X"FD",X"C4",X"FE",X"D8",X"03",X"04",X"02",X"C4",X"FE",X"31",X"00",
		X"00",X"B0",X"FF",X"50",X"00",X"50",X"00",X"60",X"FF",X"64",X"00",X"50",X"00",X"60",X"FF",X"78",
		X"00",X"00",X"00",X"B0",X"FF",X"8C",X"00",X"00",X"00",X"50",X"00",X"50",X"00",X"50",X"00",X"A0",
		X"00",X"64",X"00",X"50",X"00",X"A0",X"00",X"78",X"00",X"00",X"00",X"50",X"00",X"8C",X"00",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"B4",X"FD",X"A8",X"FE",X"6C",X"FF",X"B4",X"FD",X"58",
		X"01",X"6C",X"FF",X"4C",X"02",X"58",X"01",X"18",X"FE",X"4C",X"02",X"A8",X"FE",X"18",X"FE",X"F0",
		X"FE",X"58",X"FF",X"D0",X"FF",X"F0",X"FE",X"A8",X"00",X"D0",X"FF",X"00",X"00",X"D8",X"FF",X"44",
		X"FF",X"00",X"00",X"28",X"00",X"44",X"FF",X"B4",X"00",X"28",X"00",X"E0",X"FE",X"B4",X"00",X"D8",
		X"FF",X"E0",X"FE",X"38",X"04",X"28",X"00",X"0C",X"FE",X"10",X"04",X"28",X"00",X"E8",X"FD",X"38",
		X"04",X"D8",X"FF",X"0C",X"FE",X"10",X"04",X"D8",X"FF",X"E8",X"FD",X"25",X"DC",X"00",X"00",X"00",
		X"F0",X"FE",X"C0",X"FE",X"B0",X"FF",X"44",X"FF",X"54",X"01",X"50",X"00",X"A0",X"FF",X"48",X"FF",
		X"00",X"00",X"9C",X"FE",X"84",X"FF",X"B0",X"FF",X"00",X"FF",X"8C",X"FF",X"50",X"00",X"30",X"FF",
		X"31",X"10",X"FF",X"88",X"FF",X"C0",X"FE",X"88",X"FE",X"40",X"00",X"E8",X"FE",X"D0",X"02",X"A0",
		X"00",X"80",X"FE",X"80",X"02",X"88",X"FF",X"C0",X"FE",X"D8",X"FF",X"C0",X"FF",X"B0",X"FF",X"00",
		X"00",X"20",X"00",X"C4",X"FF",X"38",X"00",X"60",X"FF",X"38",X"FF",X"78",X"00",X"C8",X"00",X"10",
		X"FF",X"19",X"B0",X"FF",X"F4",X"FF",X"E0",X"FE",X"D8",X"01",X"70",X"00",X"50",X"FE",X"20",X"03",
		X"D4",X"FF",X"0C",X"00",X"58",X"00",X"F0",X"FF",X"F4",X"FE",X"31",X"D4",X"FE",X"B8",X"FF",X"48",
		X"FF",X"18",X"FF",X"58",X"FF",X"48",X"FF",X"18",X"FF",X"F0",X"FE",X"14",X"FF",X"D4",X"FE",X"F0",
		X"FE",X"E4",X"FE",X"A0",X"FF",X"A8",X"00",X"34",X"FF",X"28",X"00",X"0C",X"00",X"40",X"FF",X"28",
		X"00",X"FC",X"FE",X"BC",X"FE",X"A0",X"FF",X"18",X"FF",X"6C",X"FE",X"1F",X"E0",X"FC",X"E0",X"FC",
		X"C0",X"FE",X"E0",X"FC",X"20",X"03",X"C0",X"FE",X"20",X"03",X"20",X"03",X"C0",X"FE",X"20",X"03",
		X"E0",X"FC",X"C0",X"FE",X"00",X"00",X"00",X"00",X"90",X"01",X"31",X"80",X"FD",X"80",X"FD",X"C0",
		X"FE",X"80",X"FD",X"80",X"02",X"C0",X"FE",X"80",X"02",X"80",X"02",X"C0",X"FE",X"80",X"02",X"80",
		X"FD",X"C0",X"FE",X"80",X"FD",X"80",X"FD",X"D8",X"FF",X"80",X"FD",X"80",X"02",X"D8",X"FF",X"80",
		X"02",X"80",X"02",X"D8",X"FF",X"80",X"02",X"80",X"FD",X"D8",X"FF",X"9D",X"80",X"FE",X"90",X"00",
		X"00",X"00",X"80",X"FE",X"48",X"00",X"30",X"00",X"80",X"FE",X"B8",X"FF",X"30",X"00",X"80",X"FE",
		X"70",X"FF",X"00",X"00",X"80",X"FE",X"B8",X"FF",X"D0",X"FF",X"80",X"FE",X"48",X"00",X"D0",X"FF",
		X"A0",X"FF",X"20",X"01",X"00",X"00",X"A0",X"FF",X"C0",X"00",X"60",X"00",X"A0",X"FF",X"40",X"FF",
		X"60",X"00",X"A0",X"FF",X"E0",X"FE",X"00",X"00",X"A0",X"FF",X"40",X"FF",X"A0",X"FF",X"A0",X"FF",
		X"C0",X"00",X"A0",X"FF",X"80",X"04",X"00",X"00",X"00",X"00",X"70",X"05",X"00",X"00",X"00",X"00",
		X"70",X"FF",X"70",X"FF",X"58",X"FF",X"70",X"FF",X"90",X"00",X"58",X"FF",X"90",X"00",X"90",X"00",
		X"58",X"FF",X"90",X"00",X"70",X"FF",X"58",X"FF",X"D0",X"FF",X"D0",X"FF",X"A4",X"FF",X"D0",X"FF",
		X"30",X"00",X"A4",X"FF",X"30",X"00",X"30",X"00",X"AC",X"FF",X"30",X"00",X"D0",X"FF",X"AC",X"FF",
		X"A0",X"FF",X"00",X"00",X"60",X"00",X"10",X"02",X"48",X"00",X"30",X"00",X"10",X"02",X"B8",X"FF",
		X"30",X"00",X"30",X"00",X"00",X"00",X"90",X"00",X"31",X"00",X"00",X"34",X"00",X"4C",X"FF",X"24",
		X"00",X"24",X"00",X"4C",X"FF",X"34",X"00",X"00",X"00",X"4C",X"FF",X"24",X"00",X"DC",X"FF",X"4C",
		X"FF",X"00",X"00",X"CC",X"FF",X"4C",X"FF",X"DC",X"FF",X"DC",X"FF",X"4C",X"FF",X"CC",X"FF",X"00",
		X"00",X"4C",X"FF",X"DC",X"FF",X"24",X"00",X"4C",X"FF",X"31",X"00",X"00",X"64",X"00",X"38",X"FF",
		X"48",X"00",X"48",X"00",X"38",X"FF",X"64",X"00",X"00",X"00",X"38",X"FF",X"48",X"00",X"B8",X"FF",
		X"38",X"FF",X"00",X"00",X"9C",X"FF",X"38",X"FF",X"B8",X"FF",X"B8",X"FF",X"38",X"FF",X"9C",X"FF",
		X"00",X"00",X"38",X"FF",X"B8",X"FF",X"48",X"00",X"38",X"FF",X"31",X"00",X"00",X"98",X"00",X"24",
		X"FF",X"6C",X"00",X"6C",X"00",X"24",X"FF",X"98",X"00",X"00",X"00",X"24",X"FF",X"6C",X"00",X"94",
		X"FF",X"24",X"FF",X"00",X"00",X"68",X"FF",X"24",X"FF",X"94",X"FF",X"94",X"FF",X"24",X"FF",X"68",
		X"FF",X"00",X"00",X"24",X"FF",X"94",X"FF",X"6C",X"00",X"24",X"FF",X"31",X"00",X"00",X"C8",X"00",
		X"10",X"FF",X"90",X"00",X"90",X"00",X"10",X"FF",X"C8",X"00",X"00",X"00",X"10",X"FF",X"90",X"00",
		X"70",X"FF",X"10",X"FF",X"00",X"00",X"38",X"FF",X"10",X"FF",X"70",X"FF",X"70",X"FF",X"10",X"FF",
		X"38",X"FF",X"00",X"00",X"10",X"FF",X"70",X"FF",X"90",X"00",X"10",X"FF",X"31",X"00",X"00",X"FC",
		X"00",X"FC",X"FE",X"B0",X"00",X"B0",X"00",X"FC",X"FE",X"FC",X"00",X"00",X"00",X"FC",X"FE",X"B0",
		X"00",X"50",X"FF",X"FC",X"FE",X"00",X"00",X"04",X"FF",X"FC",X"FE",X"50",X"FF",X"50",X"FF",X"FC",
		X"FE",X"04",X"FF",X"00",X"00",X"FC",X"FE",X"50",X"FF",X"B0",X"00",X"FC",X"FE",X"31",X"00",X"00",
		X"2C",X"01",X"E8",X"FE",X"D4",X"00",X"D4",X"00",X"E8",X"FE",X"2C",X"01",X"00",X"00",X"E8",X"FE",
		X"D4",X"00",X"2C",X"FF",X"E8",X"FE",X"00",X"00",X"D4",X"FE",X"E8",X"FE",X"2C",X"FF",X"2C",X"FF",
		X"E8",X"FE",X"D4",X"FE",X"00",X"00",X"E8",X"FE",X"2C",X"FF",X"D4",X"00",X"E8",X"FE",X"31",X"00",
		X"00",X"60",X"01",X"D4",X"FE",X"08",X"01",X"08",X"01",X"D4",X"FE",X"60",X"01",X"00",X"00",X"D4",
		X"FE",X"08",X"01",X"F8",X"FE",X"D4",X"FE",X"00",X"00",X"A0",X"FE",X"D4",X"FE",X"F8",X"FE",X"F8",
		X"FE",X"D4",X"FE",X"A0",X"FE",X"00",X"00",X"D4",X"FE",X"F8",X"FE",X"08",X"01",X"D4",X"FE",X"31",
		X"00",X"00",X"90",X"01",X"C0",X"FE",X"1C",X"01",X"1C",X"01",X"C0",X"FE",X"90",X"01",X"00",X"00",
		X"C0",X"FE",X"1C",X"01",X"E4",X"FE",X"C0",X"FE",X"00",X"00",X"70",X"FE",X"C0",X"FE",X"E4",X"FE",
		X"E4",X"FE",X"C0",X"FE",X"70",X"FE",X"00",X"00",X"C0",X"FE",X"E4",X"FE",X"1C",X"01",X"C0",X"FE",
		X"67",X"10",X"FF",X"00",X"00",X"D8",X"FF",X"60",X"FF",X"A0",X"00",X"D8",X"FF",X"00",X"00",X"F0",
		X"00",X"D8",X"FF",X"A0",X"00",X"A0",X"00",X"D8",X"FF",X"F0",X"00",X"00",X"00",X"D8",X"FF",X"A0",
		X"00",X"60",X"FF",X"D8",X"FF",X"00",X"00",X"10",X"FF",X"D8",X"FF",X"60",X"FF",X"60",X"FF",X"D8",
		X"FF",X"40",X"FC",X"00",X"00",X"50",X"00",X"58",X"FD",X"A8",X"02",X"50",X"00",X"00",X"00",X"C0",
		X"03",X"50",X"00",X"A8",X"02",X"A8",X"02",X"50",X"00",X"C0",X"03",X"00",X"00",X"50",X"00",X"A8",
		X"02",X"58",X"FD",X"50",X"00",X"00",X"00",X"40",X"FC",X"50",X"00",X"58",X"FD",X"58",X"FD",X"50",
		X"00",X"00",X"00",X"00",X"00",X"18",X"01",X"97",X"B0",X"05",X"70",X"01",X"C0",X"FE",X"38",X"FE",
		X"28",X"02",X"C0",X"FE",X"38",X"FE",X"D8",X"FD",X"C0",X"FE",X"B0",X"05",X"90",X"FE",X"C0",X"FE",
		X"38",X"FE",X"C8",X"01",X"A4",X"FF",X"38",X"FE",X"38",X"FE",X"A4",X"FF",X"48",X"04",X"00",X"00",
		X"EC",X"FE",X"F0",X"FE",X"10",X"01",X"8C",X"FF",X"38",X"FE",X"10",X"01",X"A4",X"FF",X"38",X"FE",
		X"F0",X"FE",X"A4",X"FF",X"F0",X"FE",X"F0",X"FE",X"8C",X"FF",X"F0",X"FE",X"B8",X"00",X"2C",X"00",
		X"38",X"FE",X"B8",X"00",X"2C",X"00",X"38",X"FE",X"48",X"FF",X"2C",X"00",X"F0",X"FE",X"48",X"FF",
		X"2C",X"00",X"00",X"05",X"58",X"00",X"D4",X"FF",X"58",X"00",X"58",X"00",X"D4",X"FF",X"58",X"00",
		X"A8",X"FF",X"D4",X"FF",X"00",X"05",X"A8",X"FF",X"D4",X"FF",X"00",X"05",X"58",X"00",X"00",X"00",
		X"A8",X"FF",X"58",X"00",X"00",X"00",X"A8",X"FF",X"A8",X"FF",X"00",X"00",X"00",X"05",X"A8",X"FF",
		X"00",X"00",X"38",X"FE",X"00",X"00",X"2C",X"00",X"38",X"FE",X"00",X"00",X"14",X"01",X"88",X"FF",
		X"88",X"FF",X"14",X"00",X"C8",X"00",X"00",X"00",X"60",X"FF",X"78",X"00",X"00",X"00",X"EC",X"FF",
		X"C8",X"00",X"60",X"FF",X"60",X"FF",X"37",X"28",X"46",X"58",X"28",X"42",X"0C",X"00",X"0F",X"10",
		X"0C",X"20",X"0F",X"40",X"0C",X"18",X"00",X"28",X"01",X"30",X"00",X"38",X"01",X"40",X"0F",X"48",
		X"0C",X"50",X"00",X"58",X"01",X"60",X"0F",X"68",X"0C",X"70",X"00",X"78",X"01",X"80",X"0F",X"88",
		X"0C",X"90",X"00",X"98",X"01",X"A0",X"FF",X"17",X"80",X"1E",X"80",X"1F",X"80",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
